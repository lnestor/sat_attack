
module c5315 ( N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, 
        N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, 
        N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
        N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, 
        N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, 
        N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, 
        N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, 
        N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
        N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, 
        N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, 
        N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, 
        N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, 
        N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
        N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, 
        N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, 
        N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, 
        N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, 
        N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, 
        N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, 
        N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, 
        N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, 
        N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, 
        N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, 
        N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, 
        N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, 
        N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, 
        N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128, keyinput0, 
        keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, 
        keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, 
        keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, 
        keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, 
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, 
        keyinput31 );
  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37,
         N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79,
         N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106,
         N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136,
         N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164,
         N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197,
         N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234,
         N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273,
         N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
         N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358,
         N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422,
         N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545,
         N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583,
         N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610,
         N613, N616, N619, N625, N631, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060,
         N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357,
         N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737,
         N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716,
         N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449,
         N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476,
         N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520,
         N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
         N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706,
         N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754,
         N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123,
         N8124, N8127, N8128;
  wire   N1, N137, N141, N293, N299, N549, N592, N1137, N1141, N4278, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164;
  assign N3360 = N1;
  assign N3359 = N1;
  assign N3358 = N1;
  assign N3357 = N1;
  assign N2309 = N1;
  assign N2139 = N137;
  assign N2142 = N141;
  assign N709 = N141;
  assign N816 = N293;
  assign N3604 = N299;
  assign N2527 = N299;
  assign N2387 = N549;
  assign N1066 = N592;
  assign N1143 = N1137;
  assign N1142 = N1137;
  assign N2584 = N1141;
  assign N4275 = N4278;

  NAND2X0 U738 ( .IN1(n674), .IN2(N137), .QN(N8128) );
  MUX41X1 U739 ( .IN1(n675), .IN3(n676), .IN2(N179), .IN4(N176), .S0(n677), 
        .S1(N580), .Q(n674) );
  NAND2X0 U740 ( .IN1(n678), .IN2(N137), .QN(N8127) );
  MUX41X1 U741 ( .IN1(n675), .IN3(n676), .IN2(N179), .IN4(N176), .S0(n679), 
        .S1(N574), .Q(n678) );
  AO221X1 U742 ( .IN1(n680), .IN2(n675), .IN3(n681), .IN4(n676), .IN5(n682), 
        .Q(N8124) );
  AO22X1 U743 ( .IN1(N64), .IN2(n683), .IN3(N14), .IN4(n684), .Q(n682) );
  AO221X1 U744 ( .IN1(n685), .IN2(n675), .IN3(n686), .IN4(n676), .IN5(n687), 
        .Q(N8123) );
  AO22X1 U745 ( .IN1(n688), .IN2(N14), .IN3(n689), .IN4(N64), .Q(n687) );
  AO222X1 U746 ( .IN1(n690), .IN2(n691), .IN3(N94), .IN4(N625), .IN5(n692), 
        .IN6(n693), .Q(n676) );
  INVX0 U747 ( .INP(n694), .ZN(n693) );
  INVX0 U748 ( .INP(n695), .ZN(n690) );
  AO222X1 U749 ( .IN1(n691), .IN2(n696), .IN3(n692), .IN4(n697), .IN5(N97), 
        .IN6(N625), .Q(n675) );
  AO222X1 U750 ( .IN1(n698), .IN2(n691), .IN3(N619), .IN4(n699), .IN5(N118), 
        .IN6(N625), .Q(N8076) );
  NAND2X0 U751 ( .IN1(n697), .IN2(n700), .QN(n699) );
  XOR2X1 U752 ( .IN1(n701), .IN2(n702), .Q(n697) );
  MUX21X1 U753 ( .IN1(n703), .IN2(n704), .S(N566), .Q(n702) );
  XOR2X1 U754 ( .IN1(n705), .IN2(n706), .Q(n704) );
  XNOR3X1 U755 ( .IN1(n707), .IN2(n708), .IN3(n709), .Q(n706) );
  MUX21X1 U756 ( .IN1(n710), .IN2(n711), .S(n712), .Q(n709) );
  XOR2X1 U757 ( .IN1(n713), .IN2(n714), .Q(n712) );
  NOR2X0 U758 ( .IN1(n715), .IN2(n716), .QN(n714) );
  NOR2X0 U759 ( .IN1(N374), .IN2(n717), .QN(n713) );
  NOR2X0 U760 ( .IN1(n718), .IN2(n719), .QN(n711) );
  OR2X1 U761 ( .IN1(n719), .IN2(n718), .Q(n710) );
  XNOR3X1 U762 ( .IN1(n720), .IN2(n721), .IN3(n722), .Q(n705) );
  NAND2X0 U763 ( .IN1(n723), .IN2(n724), .QN(n722) );
  XNOR3X1 U764 ( .IN1(n719), .IN2(n725), .IN3(n726), .Q(n703) );
  XOR3X1 U765 ( .IN1(n727), .IN2(n708), .IN3(n728), .Q(n726) );
  XNOR3X1 U766 ( .IN1(n720), .IN2(n721), .IN3(n729), .Q(n728) );
  XNOR2X1 U767 ( .IN1(n730), .IN2(n731), .Q(n708) );
  XNOR3X1 U768 ( .IN1(keyinput30), .IN2(n732), .IN3(n716), .Q(n727) );
  MUX21X1 U769 ( .IN1(n733), .IN2(n734), .S(n735), .Q(n701) );
  AOI21X1 U770 ( .IN1(n736), .IN2(N566), .IN3(n737), .QN(n735) );
  XNOR2X1 U771 ( .IN1(n738), .IN2(n739), .Q(n734) );
  OA21X1 U772 ( .IN1(n740), .IN2(n741), .IN3(n742), .Q(n739) );
  XOR2X1 U773 ( .IN1(n743), .IN2(keyinput29), .Q(n742) );
  NAND2X0 U774 ( .IN1(n740), .IN2(n741), .QN(n743) );
  XNOR3X1 U775 ( .IN1(n744), .IN2(n745), .IN3(n746), .Q(n740) );
  XOR2X1 U776 ( .IN1(n747), .IN2(n748), .Q(n746) );
  XOR3X1 U777 ( .IN1(n748), .IN2(n749), .IN3(n750), .Q(n733) );
  MUX21X1 U778 ( .IN1(n751), .IN2(n752), .S(n753), .Q(n750) );
  NOR2X0 U779 ( .IN1(n752), .IN2(n738), .QN(n751) );
  XNOR3X1 U780 ( .IN1(n741), .IN2(n754), .IN3(n738), .Q(n749) );
  XNOR2X1 U781 ( .IN1(n755), .IN2(n756), .Q(n748) );
  INVX0 U782 ( .INP(n696), .ZN(n698) );
  XOR3X1 U783 ( .IN1(n757), .IN2(n758), .IN3(n759), .Q(n696) );
  XOR3X1 U784 ( .IN1(n760), .IN2(n761), .IN3(n762), .Q(n759) );
  NAND2X0 U785 ( .IN1(n763), .IN2(n764), .QN(n762) );
  XNOR2X1 U786 ( .IN1(n765), .IN2(keyinput19), .Q(n764) );
  NAND3X0 U787 ( .IN1(n766), .IN2(n767), .IN3(n768), .QN(n765) );
  MUX21X1 U788 ( .IN1(n769), .IN2(n770), .S(n768), .Q(n763) );
  XOR2X1 U789 ( .IN1(n771), .IN2(n772), .Q(n768) );
  MUX41X1 U790 ( .IN1(N251), .IN3(N248), .IN2(n773), .IN4(n774), .S0(N273), 
        .S1(n775), .Q(n772) );
  MUX41X1 U791 ( .IN1(N254), .IN3(n776), .IN2(N242), .IN4(n777), .S0(N400), 
        .S1(N265), .Q(n771) );
  OR2X1 U792 ( .IN1(n766), .IN2(n767), .Q(n770) );
  XNOR2X1 U793 ( .IN1(n766), .IN2(n767), .Q(n769) );
  XNOR2X1 U794 ( .IN1(n778), .IN2(n779), .Q(n767) );
  MUX41X1 U795 ( .IN1(N251), .IN3(N248), .IN2(n773), .IN4(n774), .S0(N257), 
        .S1(n780), .Q(n779) );
  MUX41X1 U796 ( .IN1(n776), .IN3(N254), .IN2(n777), .IN4(N242), .S0(n781), 
        .S1(N234), .Q(n778) );
  MUX41X1 U797 ( .IN1(n776), .IN3(N254), .IN2(n777), .IN4(N242), .S0(n782), 
        .S1(N281), .Q(n766) );
  MUX41X1 U798 ( .IN1(n773), .IN3(n774), .IN2(N251), .IN4(N248), .S0(N226), 
        .S1(N422), .Q(n761) );
  OA21X1 U799 ( .IN1(keyinput7), .IN2(n783), .IN3(n784), .Q(n760) );
  MUX21X1 U800 ( .IN1(n785), .IN2(n786), .S(n787), .Q(n784) );
  MUX21X1 U801 ( .IN1(N254), .IN2(N242), .S(N210), .Q(n786) );
  NAND2X0 U802 ( .IN1(keyinput7), .IN2(n788), .QN(n785) );
  MUX21X1 U803 ( .IN1(N251), .IN2(N248), .S(N210), .Q(n788) );
  AND3X1 U804 ( .IN1(N457), .IN2(N210), .IN3(N248), .Q(n783) );
  MUX41X1 U805 ( .IN1(n773), .IN3(n774), .IN2(N251), .IN4(N248), .S0(N218), 
        .S1(N468), .Q(n757) );
  AO221X1 U806 ( .IN1(N625), .IN2(n789), .IN3(n691), .IN4(n695), .IN5(n790), 
        .Q(N8075) );
  XOR2X1 U807 ( .IN1(n791), .IN2(keyinput31), .Q(n790) );
  NAND2X0 U808 ( .IN1(n694), .IN2(N619), .QN(n791) );
  XOR3X1 U809 ( .IN1(n792), .IN2(n793), .IN3(n794), .Q(n694) );
  MUX21X1 U810 ( .IN1(n795), .IN2(n796), .S(N583), .Q(n794) );
  XOR3X1 U811 ( .IN1(n797), .IN2(n798), .IN3(n799), .Q(n796) );
  MUX21X1 U812 ( .IN1(n800), .IN2(n801), .S(n802), .Q(n799) );
  NAND2X0 U813 ( .IN1(n803), .IN2(n804), .QN(n801) );
  OA21X1 U814 ( .IN1(n805), .IN2(n804), .IN3(n803), .Q(n800) );
  INVX0 U815 ( .INP(n806), .ZN(n803) );
  XOR3X1 U816 ( .IN1(n807), .IN2(n808), .IN3(n809), .Q(n798) );
  NAND3X0 U817 ( .IN1(n810), .IN2(n811), .IN3(n812), .QN(n809) );
  NAND2X0 U818 ( .IN1(n813), .IN2(n814), .QN(n810) );
  XNOR2X1 U819 ( .IN1(n815), .IN2(n816), .Q(n797) );
  XOR3X1 U820 ( .IN1(n817), .IN2(n818), .IN3(n819), .Q(n795) );
  XOR2X1 U821 ( .IN1(n820), .IN2(n821), .Q(n819) );
  OA21X1 U822 ( .IN1(n822), .IN2(n823), .IN3(n824), .Q(n821) );
  XOR2X1 U823 ( .IN1(keyinput22), .IN2(n825), .Q(n824) );
  NOR2X0 U824 ( .IN1(n816), .IN2(n802), .QN(n825) );
  INVX0 U825 ( .INP(n802), .ZN(n822) );
  AO21X1 U826 ( .IN1(n805), .IN2(n806), .IN3(n826), .Q(n802) );
  NAND2X0 U827 ( .IN1(n827), .IN2(n812), .QN(n820) );
  NOR2X0 U828 ( .IN1(n828), .IN2(n829), .QN(n812) );
  AND3X1 U829 ( .IN1(n814), .IN2(n808), .IN3(n816), .Q(n829) );
  XNOR2X1 U830 ( .IN1(n830), .IN2(keyinput18), .Q(n827) );
  XNOR2X1 U831 ( .IN1(n808), .IN2(n806), .Q(n818) );
  XNOR3X1 U832 ( .IN1(n807), .IN2(n815), .IN3(n816), .Q(n817) );
  XNOR2X1 U833 ( .IN1(n831), .IN2(n805), .Q(n807) );
  MUX21X1 U834 ( .IN1(n832), .IN2(n833), .S(n834), .Q(n793) );
  NOR2X0 U835 ( .IN1(n835), .IN2(n836), .QN(n834) );
  AND3X1 U836 ( .IN1(N583), .IN2(n813), .IN3(n837), .Q(n835) );
  INVX0 U837 ( .INP(n804), .ZN(n813) );
  XOR3X1 U838 ( .IN1(n838), .IN2(n839), .IN3(n840), .Q(n833) );
  XOR3X1 U839 ( .IN1(n841), .IN2(n839), .IN3(n842), .Q(n832) );
  OR2X1 U840 ( .IN1(n843), .IN2(n844), .Q(n842) );
  NOR2X0 U841 ( .IN1(n845), .IN2(n846), .QN(n792) );
  MUX21X1 U842 ( .IN1(n847), .IN2(n848), .S(n849), .Q(n846) );
  NOR2X0 U843 ( .IN1(n850), .IN2(n851), .QN(n848) );
  XNOR2X1 U844 ( .IN1(n851), .IN2(n852), .Q(n847) );
  XNOR3X1 U845 ( .IN1(n853), .IN2(n854), .IN3(n855), .Q(n695) );
  XOR2X1 U846 ( .IN1(n856), .IN2(n857), .Q(n855) );
  OA21X1 U847 ( .IN1(n858), .IN2(n859), .IN3(n860), .Q(n857) );
  XOR2X1 U848 ( .IN1(keyinput13), .IN2(n861), .Q(n860) );
  AND2X1 U849 ( .IN1(n859), .IN2(n858), .Q(n861) );
  MUX21X1 U850 ( .IN1(n862), .IN2(n863), .S(n864), .Q(n856) );
  AND2X1 U851 ( .IN1(n865), .IN2(n866), .Q(n863) );
  NAND2X0 U852 ( .IN1(n866), .IN2(n865), .QN(n862) );
  XNOR3X1 U853 ( .IN1(n867), .IN2(n868), .IN3(n869), .Q(n854) );
  MUX41X1 U854 ( .IN1(n776), .IN3(N254), .IN2(n777), .IN4(N242), .S0(n870), 
        .S1(N351), .Q(n869) );
  MUX41X1 U855 ( .IN1(N251), .IN3(N248), .IN2(n773), .IN4(n774), .S0(N341), 
        .S1(n871), .Q(n867) );
  MUX21X1 U856 ( .IN1(n872), .IN2(n873), .S(N514), .Q(n853) );
  XNOR2X1 U857 ( .IN1(n874), .IN2(n777), .Q(n873) );
  XNOR2X1 U858 ( .IN1(N242), .IN2(n874), .Q(n872) );
  MUX41X1 U859 ( .IN1(n776), .IN3(N254), .IN2(n777), .IN4(N242), .S0(n875), 
        .S1(N324), .Q(n874) );
  OR2X1 U860 ( .IN1(N120), .IN2(N619), .Q(n789) );
  AO221X1 U861 ( .IN1(n876), .IN2(n877), .IN3(N161), .IN4(n878), .IN5(n879), 
        .Q(N7761) );
  AO22X1 U862 ( .IN1(N191), .IN2(n880), .IN3(n881), .IN4(n882), .Q(n879) );
  AO221X1 U863 ( .IN1(n881), .IN2(n883), .IN3(n876), .IN4(n884), .IN5(n885), 
        .Q(N7760) );
  AO22X1 U864 ( .IN1(N164), .IN2(n878), .IN3(N194), .IN4(n880), .Q(n885) );
  AO221X1 U865 ( .IN1(N167), .IN2(n878), .IN3(n881), .IN4(n886), .IN5(n887), 
        .Q(N7759) );
  AO22X1 U866 ( .IN1(N197), .IN2(n880), .IN3(n876), .IN4(n888), .Q(n887) );
  AO221X1 U867 ( .IN1(n876), .IN2(n889), .IN3(N203), .IN4(n880), .IN5(n890), 
        .Q(N7758) );
  AO22X1 U868 ( .IN1(n881), .IN2(n891), .IN3(N173), .IN4(n878), .Q(n890) );
  AO221X1 U869 ( .IN1(n892), .IN2(n882), .IN3(n893), .IN4(n877), .IN5(n894), 
        .Q(N7757) );
  AO22X1 U870 ( .IN1(n895), .IN2(N161), .IN3(n896), .IN4(N191), .Q(n894) );
  AO221X1 U871 ( .IN1(n892), .IN2(n883), .IN3(n893), .IN4(n884), .IN5(n897), 
        .Q(N7756) );
  AO22X1 U872 ( .IN1(n895), .IN2(N164), .IN3(n896), .IN4(N194), .Q(n897) );
  AO221X1 U873 ( .IN1(n895), .IN2(N167), .IN3(n892), .IN4(n886), .IN5(n898), 
        .Q(N7755) );
  AO22X1 U874 ( .IN1(n896), .IN2(N197), .IN3(n893), .IN4(n888), .Q(n898) );
  AO221X1 U875 ( .IN1(n893), .IN2(n889), .IN3(n896), .IN4(N203), .IN5(n899), 
        .Q(N7754) );
  AO22X1 U876 ( .IN1(n892), .IN2(n891), .IN3(n895), .IN4(N173), .Q(n899) );
  AO221X1 U877 ( .IN1(n681), .IN2(n889), .IN3(N91), .IN4(n684), .IN5(n900), 
        .Q(N7742) );
  AO22X1 U878 ( .IN1(n680), .IN2(n891), .IN3(N40), .IN4(n683), .Q(n900) );
  AO221X1 U879 ( .IN1(N103), .IN2(n683), .IN3(n680), .IN4(n886), .IN5(n901), 
        .Q(N7741) );
  AO22X1 U880 ( .IN1(N100), .IN2(n684), .IN3(n681), .IN4(n888), .Q(n901) );
  AO221X1 U881 ( .IN1(n680), .IN2(n883), .IN3(n681), .IN4(n884), .IN5(n902), 
        .Q(N7740) );
  AO22X1 U882 ( .IN1(N49), .IN2(n683), .IN3(N46), .IN4(n684), .Q(n902) );
  AO221X1 U883 ( .IN1(n686), .IN2(n889), .IN3(N40), .IN4(n689), .IN5(n903), 
        .Q(N7739) );
  AO21X1 U884 ( .IN1(N91), .IN2(n688), .IN3(n904), .Q(n903) );
  XOR2X1 U885 ( .IN1(n905), .IN2(keyinput28), .Q(n904) );
  NAND2X0 U886 ( .IN1(n685), .IN2(n891), .QN(n905) );
  AO221X1 U887 ( .IN1(n686), .IN2(n888), .IN3(N100), .IN4(n688), .IN5(n906), 
        .Q(N7738) );
  AO21X1 U888 ( .IN1(n685), .IN2(n886), .IN3(n907), .Q(n906) );
  XOR2X1 U889 ( .IN1(n908), .IN2(keyinput2), .Q(n907) );
  NAND2X0 U890 ( .IN1(N103), .IN2(n689), .QN(n908) );
  AO221X1 U891 ( .IN1(n685), .IN2(n883), .IN3(N49), .IN4(n689), .IN5(n909), 
        .Q(N7737) );
  AO21X1 U892 ( .IN1(N46), .IN2(n688), .IN3(n910), .Q(n909) );
  XOR2X1 U893 ( .IN1(keyinput27), .IN2(n911), .Q(n910) );
  AND2X1 U894 ( .IN1(n884), .IN2(n686), .Q(n911) );
  AO221X1 U895 ( .IN1(N109), .IN2(n688), .IN3(n686), .IN4(n877), .IN5(n912), 
        .Q(N7736) );
  AO22X1 U896 ( .IN1(N106), .IN2(n689), .IN3(n685), .IN4(n882), .Q(n912) );
  AO221X1 U897 ( .IN1(n680), .IN2(n882), .IN3(N109), .IN4(n684), .IN5(n913), 
        .Q(N7735) );
  AO21X1 U898 ( .IN1(n681), .IN2(n877), .IN3(n914), .Q(n913) );
  XOR2X1 U899 ( .IN1(keyinput1), .IN2(n915), .Q(n914) );
  AND2X1 U900 ( .IN1(n683), .IN2(N106), .Q(n915) );
  INVX0 U901 ( .INP(n891), .ZN(N7707) );
  AO221X1 U902 ( .IN1(n916), .IN2(n691), .IN3(n917), .IN4(n692), .IN5(n918), 
        .Q(n891) );
  XOR2X1 U903 ( .IN1(n919), .IN2(keyinput10), .Q(n918) );
  NAND2X0 U904 ( .IN1(N113), .IN2(n920), .QN(n919) );
  INVX0 U905 ( .INP(n886), .ZN(N7706) );
  AO222X1 U906 ( .IN1(n921), .IN2(n691), .IN3(N53), .IN4(n920), .IN5(n922), 
        .IN6(n692), .Q(n886) );
  INVX0 U907 ( .INP(n883), .ZN(N7705) );
  AO222X1 U908 ( .IN1(N114), .IN2(n920), .IN3(n923), .IN4(n692), .IN5(n924), 
        .IN6(n691), .Q(n883) );
  MUX21X1 U909 ( .IN1(n925), .IN2(n926), .S(n927), .Q(n923) );
  XOR2X1 U910 ( .IN1(n745), .IN2(n928), .Q(n925) );
  INVX0 U911 ( .INP(n882), .ZN(N7704) );
  AO222X1 U912 ( .IN1(N115), .IN2(n920), .IN3(n692), .IN4(n929), .IN5(n691), 
        .IN6(n758), .Q(n882) );
  NOR2X0 U913 ( .IN1(n930), .IN2(n931), .QN(N7703) );
  OR4X1 U914 ( .IN1(n932), .IN2(N6877), .IN3(N7476), .IN4(N6716), .Q(n931) );
  INVX0 U915 ( .INP(N1140), .ZN(n932) );
  OR4X1 U916 ( .IN1(N1152), .IN2(N1155), .IN3(N2061), .IN4(N7474), .Q(n930) );
  INVX0 U917 ( .INP(n889), .ZN(N7702) );
  AO222X1 U918 ( .IN1(N112), .IN2(n920), .IN3(n933), .IN4(n692), .IN5(n864), 
        .IN6(n691), .Q(n889) );
  INVX0 U919 ( .INP(n888), .ZN(N7701) );
  AO222X1 U920 ( .IN1(N116), .IN2(n920), .IN3(n692), .IN4(n934), .IN5(n935), 
        .IN6(n691), .Q(n888) );
  INVX0 U921 ( .INP(n884), .ZN(N7700) );
  AO221X1 U922 ( .IN1(N121), .IN2(n920), .IN3(n691), .IN4(n859), .IN5(n936), 
        .Q(n884) );
  XOR2X1 U923 ( .IN1(keyinput26), .IN2(n937), .Q(n936) );
  AND2X1 U924 ( .IN1(n692), .IN2(n938), .Q(n937) );
  INVX0 U925 ( .INP(n877), .ZN(N7699) );
  AO222X1 U926 ( .IN1(n692), .IN2(n939), .IN3(N123), .IN4(n920), .IN5(n940), 
        .IN6(n691), .Q(n877) );
  XNOR2X1 U927 ( .IN1(N7432), .IN2(n941), .Q(N7698) );
  AOI21X1 U928 ( .IN1(N631), .IN2(N135), .IN3(n942), .QN(N7626) );
  INVX0 U929 ( .INP(n943), .ZN(n942) );
  MUX41X1 U930 ( .IN1(n940), .IN3(n941), .IN2(N123), .IN4(n939), .S0(N603), 
        .S1(N599), .Q(n943) );
  XOR2X1 U931 ( .IN1(n944), .IN2(N132), .Q(n941) );
  AO221X1 U932 ( .IN1(n945), .IN2(n946), .IN3(N149), .IN4(n947), .IN5(n948), 
        .Q(N7607) );
  AO22X1 U933 ( .IN1(n881), .IN2(n949), .IN3(N146), .IN4(n878), .Q(n948) );
  AO221X1 U934 ( .IN1(n945), .IN2(n950), .IN3(N155), .IN4(n947), .IN5(n951), 
        .Q(N7606) );
  AO22X1 U935 ( .IN1(n881), .IN2(n952), .IN3(N152), .IN4(n878), .Q(n951) );
  AO221X1 U936 ( .IN1(N158), .IN2(n878), .IN3(n881), .IN4(n953), .IN5(n954), 
        .Q(N7605) );
  AO22X1 U937 ( .IN1(N188), .IN2(n947), .IN3(n945), .IN4(n955), .Q(n954) );
  AO221X1 U938 ( .IN1(N200), .IN2(n880), .IN3(n876), .IN4(n956), .IN5(n957), 
        .Q(N7604) );
  AO21X1 U939 ( .IN1(n878), .IN2(N170), .IN3(n958), .Q(n957) );
  INVX0 U940 ( .INP(n959), .ZN(n958) );
  MUX21X1 U941 ( .IN1(n960), .IN2(n961), .S(keyinput25), .Q(n959) );
  NAND2X0 U942 ( .IN1(N137), .IN2(n962), .QN(n961) );
  NAND3X0 U943 ( .IN1(n963), .IN2(n964), .IN3(N577), .QN(n962) );
  NAND2X0 U944 ( .IN1(n881), .IN2(n963), .QN(n960) );
  AND2X1 U945 ( .IN1(n965), .IN2(n966), .Q(n876) );
  AND2X1 U946 ( .IN1(n967), .IN2(n965), .Q(n880) );
  XNOR2X1 U947 ( .IN1(N577), .IN2(keyinput6), .Q(n965) );
  AO221X1 U948 ( .IN1(n893), .IN2(n946), .IN3(N149), .IN4(n896), .IN5(n968), 
        .Q(N7603) );
  AO22X1 U949 ( .IN1(n892), .IN2(n949), .IN3(N146), .IN4(n895), .Q(n968) );
  AO221X1 U950 ( .IN1(n893), .IN2(n950), .IN3(N155), .IN4(n896), .IN5(n969), 
        .Q(N7602) );
  AO22X1 U951 ( .IN1(n892), .IN2(n952), .IN3(N152), .IN4(n895), .Q(n969) );
  AO221X1 U952 ( .IN1(N158), .IN2(n895), .IN3(n892), .IN4(n953), .IN5(n970), 
        .Q(N7601) );
  AO22X1 U953 ( .IN1(N188), .IN2(n896), .IN3(n893), .IN4(n955), .Q(n970) );
  AO221X1 U954 ( .IN1(n893), .IN2(n956), .IN3(N200), .IN4(n896), .IN5(n971), 
        .Q(N7600) );
  AO22X1 U955 ( .IN1(n892), .IN2(n963), .IN3(N170), .IN4(n895), .Q(n971) );
  AO221X1 U956 ( .IN1(n680), .IN2(n953), .IN3(n681), .IN4(n955), .IN5(n972), 
        .Q(N7522) );
  AO22X1 U957 ( .IN1(N70), .IN2(n683), .IN3(N67), .IN4(n684), .Q(n972) );
  AO221X1 U958 ( .IN1(n680), .IN2(n952), .IN3(n681), .IN4(n950), .IN5(n973), 
        .Q(N7521) );
  AO22X1 U959 ( .IN1(N17), .IN2(n683), .IN3(N73), .IN4(n684), .Q(n973) );
  AO221X1 U960 ( .IN1(n680), .IN2(n949), .IN3(N76), .IN4(n684), .IN5(n974), 
        .Q(N7520) );
  AO21X1 U961 ( .IN1(n681), .IN2(n946), .IN3(n975), .Q(n974) );
  XOR2X1 U962 ( .IN1(n976), .IN2(keyinput4), .Q(n975) );
  NAND2X0 U963 ( .IN1(N20), .IN2(n683), .QN(n976) );
  AO221X1 U964 ( .IN1(n680), .IN2(n963), .IN3(N43), .IN4(n684), .IN5(n977), 
        .Q(N7519) );
  AO21X1 U965 ( .IN1(n681), .IN2(n956), .IN3(n978), .Q(n977) );
  XOR2X1 U966 ( .IN1(keyinput3), .IN2(n979), .Q(n978) );
  AND2X1 U967 ( .IN1(n683), .IN2(N37), .Q(n979) );
  AO221X1 U968 ( .IN1(n685), .IN2(n953), .IN3(n686), .IN4(n955), .IN5(n980), 
        .Q(N7518) );
  AO22X1 U969 ( .IN1(N67), .IN2(n688), .IN3(N70), .IN4(n689), .Q(n980) );
  AO221X1 U970 ( .IN1(n686), .IN2(n950), .IN3(N17), .IN4(n689), .IN5(n981), 
        .Q(N7517) );
  AO22X1 U971 ( .IN1(n685), .IN2(n952), .IN3(N73), .IN4(n688), .Q(n981) );
  AO221X1 U972 ( .IN1(n685), .IN2(n949), .IN3(n686), .IN4(n946), .IN5(n982), 
        .Q(N7516) );
  AO22X1 U973 ( .IN1(N76), .IN2(n688), .IN3(N20), .IN4(n689), .Q(n982) );
  AO221X1 U974 ( .IN1(n685), .IN2(n963), .IN3(n686), .IN4(n956), .IN5(n983), 
        .Q(N7515) );
  AO22X1 U975 ( .IN1(N43), .IN2(n688), .IN3(N37), .IN4(n689), .Q(n983) );
  AO221X1 U976 ( .IN1(N185), .IN2(n878), .IN3(n881), .IN4(n984), .IN5(n985), 
        .Q(N7511) );
  AO22X1 U977 ( .IN1(N182), .IN2(n947), .IN3(n945), .IN4(n986), .Q(n985) );
  AND2X1 U978 ( .IN1(n966), .IN2(n677), .Q(n945) );
  AND2X1 U979 ( .IN1(n967), .IN2(n677), .Q(n947) );
  INVX0 U980 ( .INP(N577), .ZN(n677) );
  AND2X1 U981 ( .IN1(n966), .IN2(N577), .Q(n881) );
  AND2X1 U982 ( .IN1(N137), .IN2(n964), .Q(n966) );
  INVX0 U983 ( .INP(N580), .ZN(n964) );
  AND2X1 U984 ( .IN1(n967), .IN2(N577), .Q(n878) );
  AND2X1 U985 ( .IN1(N137), .IN2(N580), .Q(n967) );
  AO221X1 U986 ( .IN1(N185), .IN2(n895), .IN3(n892), .IN4(n984), .IN5(n987), 
        .Q(N7506) );
  AO22X1 U987 ( .IN1(N182), .IN2(n896), .IN3(n893), .IN4(n986), .Q(n987) );
  AND3X1 U988 ( .IN1(n679), .IN2(n988), .IN3(N137), .Q(n893) );
  AND3X1 U989 ( .IN1(N137), .IN2(n679), .IN3(N574), .Q(n896) );
  INVX0 U990 ( .INP(N571), .ZN(n679) );
  AND3X1 U991 ( .IN1(N137), .IN2(n988), .IN3(N571), .Q(n892) );
  INVX0 U992 ( .INP(N574), .ZN(n988) );
  AND3X1 U993 ( .IN1(N571), .IN2(N137), .IN3(N574), .Q(n895) );
  NOR4X0 U994 ( .IN1(n989), .IN2(n990), .IN3(n991), .IN4(n992), .QN(N7504) );
  OR3X1 U995 ( .IN1(n933), .IN2(n938), .IN3(n993), .Q(n990) );
  OA21X1 U996 ( .IN1(n840), .IN2(n994), .IN3(n995), .Q(n938) );
  MUX21X1 U997 ( .IN1(n996), .IN2(n843), .S(n839), .Q(n995) );
  AOI21X1 U998 ( .IN1(n843), .IN2(n994), .IN3(n997), .QN(n996) );
  NAND2X0 U999 ( .IN1(n998), .IN2(n999), .QN(n843) );
  NAND2X0 U1000 ( .IN1(n998), .IN2(n997), .QN(n840) );
  INVX0 U1001 ( .INP(n1000), .ZN(n998) );
  XOR2X1 U1002 ( .IN1(n849), .IN2(n994), .Q(n933) );
  OR4X1 U1003 ( .IN1(n934), .IN2(n1001), .IN3(n1002), .IN4(n939), .Q(n989) );
  INVX0 U1004 ( .INP(N7432), .ZN(n939) );
  INVX0 U1005 ( .INP(n1003), .ZN(n934) );
  MUX21X1 U1006 ( .IN1(n1004), .IN2(n1005), .S(n994), .Q(n1003) );
  INVX0 U1007 ( .INP(n1006), .ZN(n994) );
  XNOR2X1 U1008 ( .IN1(n841), .IN2(n1007), .Q(n1005) );
  NOR2X0 U1009 ( .IN1(n1008), .IN2(N490), .QN(n841) );
  OA21X1 U1010 ( .IN1(n838), .IN2(n1007), .IN3(n1009), .Q(n1004) );
  XOR2X1 U1011 ( .IN1(n1010), .IN2(keyinput21), .Q(n1009) );
  NAND2X0 U1012 ( .IN1(n838), .IN2(n1007), .QN(n1010) );
  INVX0 U1013 ( .INP(n851), .ZN(n1007) );
  NOR4X0 U1014 ( .IN1(n1011), .IN2(n1012), .IN3(n917), .IN4(n1013), .QN(N7503)
         );
  XOR2X1 U1015 ( .IN1(n927), .IN2(n756), .Q(n917) );
  OR3X1 U1016 ( .IN1(n926), .IN2(n1014), .IN3(n922), .Q(n1012) );
  MUX21X1 U1017 ( .IN1(n1015), .IN2(n1016), .S(n755), .Q(n922) );
  AOI21X1 U1018 ( .IN1(n927), .IN2(n754), .IN3(n744), .QN(n1016) );
  OA21X1 U1019 ( .IN1(n744), .IN2(n927), .IN3(n754), .Q(n1015) );
  INVX0 U1020 ( .INP(n1017), .ZN(n754) );
  XNOR2X1 U1021 ( .IN1(n928), .IN2(n753), .Q(n926) );
  NOR2X0 U1022 ( .IN1(n745), .IN2(n1018), .QN(n753) );
  OR4X1 U1023 ( .IN1(n929), .IN2(n1019), .IN3(n1020), .IN4(n1021), .Q(n1011)
         );
  INVX0 U1024 ( .INP(n1022), .ZN(n929) );
  MUX21X1 U1025 ( .IN1(n1023), .IN2(n1024), .S(n927), .Q(n1022) );
  AO21X1 U1026 ( .IN1(N4), .IN2(n736), .IN3(n737), .Q(n927) );
  XNOR2X1 U1027 ( .IN1(n741), .IN2(n1025), .Q(n1024) );
  AOI21X1 U1028 ( .IN1(n928), .IN2(n1018), .IN3(n1026), .QN(n1025) );
  INVX0 U1029 ( .INP(n1027), .ZN(n1018) );
  XNOR3X1 U1030 ( .IN1(keyinput20), .IN2(n1028), .IN3(n1026), .Q(n1023) );
  AO21X1 U1031 ( .IN1(n1029), .IN2(n1030), .IN3(n1031), .Q(N7474) );
  XOR2X1 U1032 ( .IN1(n1032), .IN2(keyinput23), .Q(n1031) );
  OR2X1 U1033 ( .IN1(n1030), .IN2(n1029), .Q(n1032) );
  XNOR3X1 U1034 ( .IN1(n1008), .IN2(n839), .IN3(n1033), .Q(n1030) );
  XNOR2X1 U1035 ( .IN1(n944), .IN2(n1034), .Q(n1033) );
  XNOR3X1 U1036 ( .IN1(n1035), .IN2(n1036), .IN3(n1037), .Q(n1029) );
  XNOR3X1 U1037 ( .IN1(n1038), .IN2(n1039), .IN3(n1040), .Q(n1037) );
  MUX21X1 U1038 ( .IN1(n1041), .IN2(n1042), .S(N332), .Q(n1035) );
  XNOR2X1 U1039 ( .IN1(n823), .IN2(N372), .Q(n1042) );
  XNOR2X1 U1040 ( .IN1(n823), .IN2(N369), .Q(n1041) );
  INVX0 U1041 ( .INP(n953), .ZN(N7473) );
  AO222X1 U1042 ( .IN1(n1043), .IN2(n691), .IN3(N126), .IN4(n920), .IN5(n1014), 
        .IN6(n692), .Q(n953) );
  AOI21X1 U1043 ( .IN1(N4), .IN2(n718), .IN3(n1044), .QN(n1014) );
  MUX21X1 U1044 ( .IN1(n1045), .IN2(n1046), .S(n1047), .Q(n1044) );
  OA21X1 U1045 ( .IN1(n707), .IN2(n1048), .IN3(n730), .Q(n1046) );
  INVX0 U1046 ( .INP(n952), .ZN(N7472) );
  AO222X1 U1047 ( .IN1(n1049), .IN2(n691), .IN3(N127), .IN4(n920), .IN5(n1021), 
        .IN6(n692), .Q(n952) );
  XOR2X1 U1048 ( .IN1(n1050), .IN2(n721), .Q(n1021) );
  INVX0 U1049 ( .INP(n949), .ZN(N7471) );
  AO222X1 U1050 ( .IN1(N128), .IN2(n920), .IN3(n1013), .IN4(n692), .IN5(n1051), 
        .IN6(n691), .Q(n949) );
  XNOR2X1 U1051 ( .IN1(n1052), .IN2(n1053), .Q(n1013) );
  INVX0 U1052 ( .INP(n963), .ZN(N7470) );
  AO222X1 U1053 ( .IN1(N122), .IN2(n920), .IN3(n1020), .IN4(n692), .IN5(n1054), 
        .IN6(n691), .Q(n963) );
  XOR2X1 U1054 ( .IN1(n1055), .IN2(n1056), .Q(n1020) );
  OA21X1 U1055 ( .IN1(n1052), .IN2(n720), .IN3(n1057), .Q(n1056) );
  AOI21X1 U1056 ( .IN1(n721), .IN2(n1050), .IN3(n1058), .QN(n1052) );
  AO21X1 U1057 ( .IN1(N4), .IN2(n718), .IN3(n719), .Q(n1050) );
  AO221X1 U1058 ( .IN1(n680), .IN2(n984), .IN3(n681), .IN4(n986), .IN5(n1059), 
        .Q(N7469) );
  AO22X1 U1059 ( .IN1(N61), .IN2(n683), .IN3(N11), .IN4(n684), .Q(n1059) );
  AND2X1 U1060 ( .IN1(N616), .IN2(n1060), .Q(n684) );
  AND2X1 U1061 ( .IN1(N616), .IN2(N613), .Q(n683) );
  NOR2X0 U1062 ( .IN1(N613), .IN2(N616), .QN(n681) );
  NOR2X0 U1063 ( .IN1(n1060), .IN2(N616), .QN(n680) );
  INVX0 U1064 ( .INP(N613), .ZN(n1060) );
  INVX0 U1065 ( .INP(n950), .ZN(N7467) );
  AO222X1 U1066 ( .IN1(N119), .IN2(n920), .IN3(n991), .IN4(n692), .IN5(n1061), 
        .IN6(n691), .Q(n950) );
  XOR2X1 U1067 ( .IN1(n1062), .IN2(n805), .Q(n991) );
  INVX0 U1068 ( .INP(n946), .ZN(N7466) );
  AO222X1 U1069 ( .IN1(n993), .IN2(n692), .IN3(n691), .IN4(n1063), .IN5(N130), 
        .IN6(n920), .Q(n946) );
  XOR2X1 U1070 ( .IN1(n1064), .IN2(n831), .Q(n993) );
  INVX0 U1071 ( .INP(n956), .ZN(N7465) );
  AO222X1 U1072 ( .IN1(N52), .IN2(n920), .IN3(n1002), .IN4(n692), .IN5(n1065), 
        .IN6(n691), .Q(n956) );
  XNOR2X1 U1073 ( .IN1(n815), .IN2(n1066), .Q(n1002) );
  OA21X1 U1074 ( .IN1(n1064), .IN2(n831), .IN3(n1067), .Q(n1066) );
  INVX0 U1075 ( .INP(n1068), .ZN(n831) );
  AOI21X1 U1076 ( .IN1(n805), .IN2(n1062), .IN3(n826), .QN(n1064) );
  AO21X1 U1077 ( .IN1(n1069), .IN2(n1070), .IN3(n1071), .Q(n1062) );
  AO221X1 U1078 ( .IN1(n685), .IN2(n984), .IN3(n686), .IN4(n986), .IN5(n1072), 
        .Q(N7449) );
  AO22X1 U1079 ( .IN1(N11), .IN2(n688), .IN3(N61), .IN4(n689), .Q(n1072) );
  AND2X1 U1080 ( .IN1(N607), .IN2(N610), .Q(n689) );
  AND2X1 U1081 ( .IN1(N607), .IN2(n1073), .Q(n688) );
  NOR2X0 U1082 ( .IN1(N607), .IN2(N610), .QN(n686) );
  NOR2X0 U1083 ( .IN1(n1073), .IN2(N607), .QN(n685) );
  INVX0 U1084 ( .INP(N610), .ZN(n1073) );
  XOR2X1 U1085 ( .IN1(n944), .IN2(n1074), .Q(N7432) );
  OA21X1 U1086 ( .IN1(n844), .IN2(n1006), .IN3(n1075), .Q(n1074) );
  OA21X1 U1087 ( .IN1(n1076), .IN2(n1077), .IN3(n1078), .Q(n1006) );
  INVX0 U1088 ( .INP(n1079), .ZN(n1078) );
  NOR2X0 U1089 ( .IN1(n997), .IN2(n1080), .QN(n844) );
  INVX0 U1090 ( .INP(n984), .ZN(N7365) );
  AO222X1 U1091 ( .IN1(N117), .IN2(n920), .IN3(n692), .IN4(n1019), .IN5(n1081), 
        .IN6(n691), .Q(n984) );
  XNOR2X1 U1092 ( .IN1(n725), .IN2(n1048), .Q(n1019) );
  INVX0 U1093 ( .INP(N4), .ZN(n1048) );
  INVX0 U1094 ( .INP(n955), .ZN(N7363) );
  AO222X1 U1095 ( .IN1(N129), .IN2(n920), .IN3(n992), .IN4(n692), .IN5(n1082), 
        .IN6(n691), .Q(n955) );
  XOR2X1 U1096 ( .IN1(n1070), .IN2(n1069), .Q(n992) );
  INVX0 U1097 ( .INP(n986), .ZN(N7015) );
  AO222X1 U1098 ( .IN1(N131), .IN2(n920), .IN3(n692), .IN4(n1001), .IN5(n691), 
        .IN6(n868), .Q(n986) );
  NOR2X0 U1099 ( .IN1(N625), .IN2(N619), .QN(n691) );
  OAI21X1 U1100 ( .IN1(n1076), .IN2(n823), .IN3(n1070), .QN(n1001) );
  NAND2X0 U1101 ( .IN1(n823), .IN2(n1076), .QN(n1070) );
  INVX0 U1102 ( .INP(N54), .ZN(n1076) );
  AND2X1 U1103 ( .IN1(N619), .IN2(n700), .Q(n692) );
  NOR2X0 U1104 ( .IN1(n700), .IN2(N619), .QN(n920) );
  INVX0 U1105 ( .INP(N625), .ZN(n700) );
  AO221X1 U1106 ( .IN1(n845), .IN2(n836), .IN3(n850), .IN4(n997), .IN5(n1083), 
        .Q(N6927) );
  INVX0 U1107 ( .INP(n1075), .ZN(n997) );
  AO21X1 U1108 ( .IN1(n837), .IN2(n806), .IN3(n1084), .Q(n836) );
  AO21X1 U1109 ( .IN1(n816), .IN2(n808), .IN3(n1071), .Q(n806) );
  AO221X1 U1110 ( .IN1(n1085), .IN2(n1086), .IN3(n1028), .IN4(n1026), .IN5(
        n1087), .Q(N6926) );
  AO21X1 U1111 ( .IN1(n928), .IN2(n745), .IN3(n752), .Q(n1026) );
  AND2X1 U1112 ( .IN1(n737), .IN2(n928), .Q(n1085) );
  NAND3X0 U1113 ( .IN1(n944), .IN2(n1088), .IN3(n1075), .QN(N6925) );
  NOR2X0 U1114 ( .IN1(n1000), .IN2(n839), .QN(n1075) );
  AO22X1 U1115 ( .IN1(N479), .IN2(n1034), .IN3(n838), .IN4(n851), .Q(n1000) );
  AND2X1 U1116 ( .IN1(N490), .IN2(n1008), .Q(n838) );
  NAND2X0 U1117 ( .IN1(n1080), .IN2(n1079), .QN(n1088) );
  AO221X1 U1118 ( .IN1(n1089), .IN2(n1069), .IN3(n830), .IN4(n815), .IN5(n1084), .Q(n1079) );
  AO22X1 U1119 ( .IN1(N503), .IN2(n1036), .IN3(n815), .IN4(n828), .Q(n1084) );
  AO21X1 U1120 ( .IN1(n826), .IN2(n1068), .IN3(n1090), .Q(n828) );
  INVX0 U1121 ( .INP(n1067), .ZN(n1090) );
  INVX0 U1122 ( .INP(n811), .ZN(n830) );
  NAND2X0 U1123 ( .IN1(n814), .IN2(n1071), .QN(n811) );
  NOR2X0 U1124 ( .IN1(n1091), .IN2(n823), .QN(n1089) );
  INVX0 U1125 ( .INP(n999), .ZN(n1080) );
  AO221X1 U1126 ( .IN1(n1092), .IN2(n1086), .IN3(n1028), .IN4(n747), .IN5(
        n1087), .Q(N6924) );
  AO21X1 U1127 ( .IN1(n745), .IN2(n738), .IN3(n752), .Q(n747) );
  NOR2X0 U1128 ( .IN1(n787), .IN2(n1093), .QN(n752) );
  AO22X1 U1129 ( .IN1(N468), .IN2(n1094), .IN3(n744), .IN4(n755), .Q(n745) );
  INVX0 U1130 ( .INP(n741), .ZN(n1028) );
  AND2X1 U1131 ( .IN1(n737), .IN2(n738), .Q(n1092) );
  AO22X1 U1132 ( .IN1(N435), .IN2(n1095), .IN3(n731), .IN4(n729), .Q(n737) );
  INVX0 U1133 ( .INP(n723), .ZN(n729) );
  OA21X1 U1134 ( .IN1(n720), .IN2(n1096), .IN3(n1057), .Q(n723) );
  NAND2X0 U1135 ( .IN1(N389), .IN2(n1097), .QN(n1057) );
  INVX0 U1136 ( .INP(n716), .ZN(n1096) );
  AO21X1 U1137 ( .IN1(n721), .IN2(n719), .IN3(n1058), .Q(n716) );
  AND2X1 U1138 ( .IN1(N400), .IN2(n1098), .Q(n1058) );
  AO22X1 U1139 ( .IN1(N411), .IN2(n1099), .IN3(n732), .IN4(n1045), .Q(n719) );
  INVX0 U1140 ( .INP(n1047), .ZN(n732) );
  NAND2X0 U1141 ( .IN1(N374), .IN2(n717), .QN(n1047) );
  INVX0 U1142 ( .INP(n1053), .ZN(n720) );
  XNOR3X1 U1143 ( .IN1(n1100), .IN2(n1101), .IN3(N206), .Q(N6877) );
  XOR3X1 U1144 ( .IN1(N226), .IN2(N218), .IN3(N210), .Q(n1101) );
  OA21X1 U1145 ( .IN1(n1102), .IN2(n1103), .IN3(n1104), .Q(n1100) );
  XOR2X1 U1146 ( .IN1(keyinput17), .IN2(n1105), .Q(n1104) );
  NOR2X0 U1147 ( .IN1(n1106), .IN2(n1107), .QN(n1105) );
  XNOR2X1 U1148 ( .IN1(n1108), .IN2(n1109), .Q(n1106) );
  XNOR2X1 U1149 ( .IN1(n1109), .IN2(n1110), .Q(n1103) );
  INVX0 U1150 ( .INP(n1108), .ZN(n1110) );
  XOR2X1 U1151 ( .IN1(N289), .IN2(N281), .Q(n1108) );
  XOR2X1 U1152 ( .IN1(N234), .IN2(N257), .Q(n1109) );
  INVX0 U1153 ( .INP(n1107), .ZN(n1102) );
  XOR2X1 U1154 ( .IN1(N265), .IN2(N273), .Q(n1107) );
  XNOR3X1 U1155 ( .IN1(n1111), .IN2(n1112), .IN3(n1113), .Q(N6716) );
  XNOR2X1 U1156 ( .IN1(N293), .IN2(n1114), .Q(n1113) );
  OA21X1 U1157 ( .IN1(N308), .IN2(n1115), .IN3(n1116), .Q(n1114) );
  XOR2X1 U1158 ( .IN1(n1117), .IN2(keyinput8), .Q(n1116) );
  NAND2X0 U1159 ( .IN1(N308), .IN2(n1115), .QN(n1117) );
  INVX0 U1160 ( .INP(N316), .ZN(n1115) );
  XOR3X1 U1161 ( .IN1(N351), .IN2(N341), .IN3(n1118), .Q(n1112) );
  XOR2X1 U1162 ( .IN1(N369), .IN2(N361), .Q(n1118) );
  XOR2X1 U1163 ( .IN1(N324), .IN2(N302), .Q(n1111) );
  AND3X1 U1164 ( .IN1(n1086), .IN2(n736), .IN3(n928), .Q(N6648) );
  XOR2X1 U1165 ( .IN1(N457), .IN2(n1119), .Q(n928) );
  NOR4X0 U1166 ( .IN1(n804), .IN2(n1091), .IN3(n1120), .IN4(n839), .QN(N6646)
         );
  INVX0 U1167 ( .INP(n845), .ZN(n1120) );
  NOR2X0 U1168 ( .IN1(n999), .IN2(n852), .QN(n845) );
  INVX0 U1169 ( .INP(n850), .ZN(n852) );
  XOR2X1 U1170 ( .IN1(n944), .IN2(keyinput12), .Q(n850) );
  INVX0 U1171 ( .INP(n1083), .ZN(n944) );
  NAND2X0 U1172 ( .IN1(n823), .IN2(n808), .QN(n804) );
  AO22X1 U1173 ( .IN1(N534), .IN2(n1121), .IN3(n1122), .IN4(n1040), .Q(n808)
         );
  NOR2X0 U1174 ( .IN1(keyinput5), .IN2(n1071), .QN(n1122) );
  NAND2X0 U1175 ( .IN1(n1071), .IN2(n1123), .QN(n1121) );
  INVX0 U1176 ( .INP(keyinput5), .ZN(n1123) );
  NOR4X0 U1177 ( .IN1(n1083), .IN2(n999), .IN3(n1077), .IN4(n839), .QN(N6643)
         );
  MUX21X1 U1178 ( .IN1(N302), .IN2(N307), .S(N332), .Q(n839) );
  NAND3X0 U1179 ( .IN1(n837), .IN2(n823), .IN3(n1069), .QN(n1077) );
  AOI21X1 U1180 ( .IN1(n1124), .IN2(n870), .IN3(n1071), .QN(n1069) );
  NOR2X0 U1181 ( .IN1(n1124), .IN2(n870), .QN(n1071) );
  INVX0 U1182 ( .INP(n1040), .ZN(n1124) );
  MUX21X1 U1183 ( .IN1(N351), .IN2(N358), .S(N332), .Q(n1040) );
  INVX0 U1184 ( .INP(n816), .ZN(n823) );
  MUX21X1 U1185 ( .IN1(N361), .IN2(N366), .S(N332), .Q(n816) );
  INVX0 U1186 ( .INP(n1091), .ZN(n837) );
  NAND2X0 U1187 ( .IN1(n814), .IN2(n815), .QN(n1091) );
  XOR2X1 U1188 ( .IN1(N503), .IN2(n1036), .Q(n815) );
  MUX21X1 U1189 ( .IN1(N324), .IN2(N331), .S(N332), .Q(n1036) );
  AND2X1 U1190 ( .IN1(n805), .IN2(n1068), .Q(n814) );
  OA21X1 U1191 ( .IN1(n1038), .IN2(N514), .IN3(n1067), .Q(n1068) );
  NAND2X0 U1192 ( .IN1(N514), .IN2(n1038), .QN(n1067) );
  NAND2X0 U1193 ( .IN1(N332), .IN2(N1144), .QN(n1038) );
  AOI21X1 U1194 ( .IN1(n1125), .IN2(n871), .IN3(n826), .QN(n805) );
  NOR2X0 U1195 ( .IN1(n871), .IN2(n1125), .QN(n826) );
  INVX0 U1196 ( .INP(n1039), .ZN(n1125) );
  MUX21X1 U1197 ( .IN1(N341), .IN2(N348), .S(N332), .Q(n1039) );
  NAND2X0 U1198 ( .IN1(n849), .IN2(n851), .QN(n999) );
  XOR2X1 U1199 ( .IN1(N479), .IN2(n1034), .Q(n851) );
  MUX21X1 U1200 ( .IN1(N308), .IN2(N315), .S(N332), .Q(n1034) );
  XOR2X1 U1201 ( .IN1(N490), .IN2(n1008), .Q(n849) );
  MUX21X1 U1202 ( .IN1(N316), .IN2(N323), .S(N332), .Q(n1008) );
  MUX21X1 U1203 ( .IN1(N293), .IN2(N299), .S(N332), .Q(n1083) );
  AND3X1 U1204 ( .IN1(n1086), .IN2(n738), .IN3(n736), .Q(N6641) );
  NOR2X0 U1205 ( .IN1(n724), .IN2(n1055), .QN(n736) );
  INVX0 U1206 ( .INP(n731), .ZN(n1055) );
  XOR2X1 U1207 ( .IN1(N435), .IN2(n1095), .Q(n731) );
  NAND2X0 U1208 ( .IN1(n715), .IN2(n1053), .QN(n724) );
  XOR2X1 U1209 ( .IN1(N389), .IN2(n1097), .Q(n1053) );
  AND2X1 U1210 ( .IN1(n718), .IN2(n721), .Q(n715) );
  XOR2X1 U1211 ( .IN1(N400), .IN2(n1098), .Q(n721) );
  NOR2X0 U1212 ( .IN1(n707), .IN2(n730), .QN(n718) );
  INVX0 U1213 ( .INP(n1045), .ZN(n730) );
  XOR2X1 U1214 ( .IN1(N411), .IN2(n1099), .Q(n1045) );
  INVX0 U1215 ( .INP(n725), .ZN(n707) );
  XOR2X1 U1216 ( .IN1(N374), .IN2(n717), .Q(n725) );
  AO21X1 U1217 ( .IN1(n1119), .IN2(n787), .IN3(n1126), .Q(n738) );
  XOR2X1 U1218 ( .IN1(n1127), .IN2(keyinput15), .Q(n1126) );
  NAND2X0 U1219 ( .IN1(N457), .IN2(n1093), .QN(n1127) );
  NOR2X0 U1220 ( .IN1(n1027), .IN2(n741), .QN(n1086) );
  AO21X1 U1221 ( .IN1(n1128), .IN2(n1129), .IN3(n1087), .Q(n741) );
  NOR2X0 U1222 ( .IN1(n1129), .IN2(n1128), .QN(n1087) );
  INVX0 U1223 ( .INP(N446), .ZN(n1129) );
  NAND2X0 U1224 ( .IN1(n756), .IN2(n755), .QN(n1027) );
  XOR2X1 U1225 ( .IN1(n1094), .IN2(N468), .Q(n755) );
  NOR2X0 U1226 ( .IN1(n744), .IN2(n1017), .QN(n756) );
  NOR2X0 U1227 ( .IN1(n1130), .IN2(N422), .QN(n1017) );
  AND2X1 U1228 ( .IN1(N422), .IN2(n1130), .Q(n744) );
  NOR4X0 U1229 ( .IN1(n1131), .IN2(n1132), .IN3(n916), .IN4(n1051), .QN(N5388)
         );
  MUX41X1 U1230 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N257), 
        .S1(n780), .Q(n1051) );
  INVX0 U1231 ( .INP(N389), .ZN(n780) );
  MUX41X1 U1232 ( .IN1(n1133), .IN3(n1134), .IN2(N597), .IN4(N598), .S0(N226), 
        .S1(N422), .Q(n916) );
  OR3X1 U1233 ( .IN1(n924), .IN2(n758), .IN3(n921), .Q(n1132) );
  MUX41X1 U1234 ( .IN1(n1133), .IN3(n1134), .IN2(N597), .IN4(N598), .S0(N218), 
        .S1(N468), .Q(n921) );
  MUX41X1 U1235 ( .IN1(N254), .IN3(n776), .IN2(N242), .IN4(n777), .S0(N446), 
        .S1(N206), .Q(n758) );
  MUX41X1 U1236 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N210), 
        .S1(n787), .Q(n924) );
  INVX0 U1237 ( .INP(N457), .ZN(n787) );
  OR4X1 U1238 ( .IN1(n1081), .IN2(n1054), .IN3(n1043), .IN4(n1049), .Q(n1131)
         );
  MUX41X1 U1239 ( .IN1(n1133), .IN3(n1134), .IN2(N597), .IN4(N598), .S0(N265), 
        .S1(N400), .Q(n1049) );
  MUX41X1 U1240 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N273), 
        .S1(n775), .Q(n1043) );
  INVX0 U1241 ( .INP(N411), .ZN(n775) );
  MUX41X1 U1242 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N234), 
        .S1(n781), .Q(n1054) );
  INVX0 U1243 ( .INP(N435), .ZN(n781) );
  MUX41X1 U1244 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N281), 
        .S1(n782), .Q(n1081) );
  INVX0 U1245 ( .INP(N374), .ZN(n782) );
  NOR4X0 U1246 ( .IN1(n1135), .IN2(n1136), .IN3(n1061), .IN4(n1065), .QN(N5240) );
  MUX41X1 U1247 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N324), 
        .S1(n875), .Q(n1065) );
  INVX0 U1248 ( .INP(N503), .ZN(n875) );
  MUX41X1 U1249 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N341), 
        .S1(n871), .Q(n1061) );
  INVX0 U1250 ( .INP(N523), .ZN(n871) );
  OR3X1 U1251 ( .IN1(n864), .IN2(n935), .IN3(n940), .Q(n1136) );
  INVX0 U1252 ( .INP(n858), .ZN(n940) );
  MUX21X1 U1253 ( .IN1(n773), .IN2(n774), .S(N293), .Q(n858) );
  AND2X1 U1254 ( .IN1(n1137), .IN2(n866), .Q(n935) );
  NAND2X0 U1255 ( .IN1(n1138), .IN2(n1139), .QN(n866) );
  INVX0 U1256 ( .INP(N479), .ZN(n1139) );
  MUX21X1 U1257 ( .IN1(n773), .IN2(n774), .S(N308), .Q(n1138) );
  INVX0 U1258 ( .INP(N242), .ZN(n774) );
  INVX0 U1259 ( .INP(N254), .ZN(n773) );
  XOR2X1 U1260 ( .IN1(n865), .IN2(keyinput11), .Q(n1137) );
  NAND2X0 U1261 ( .IN1(n1140), .IN2(N479), .QN(n865) );
  MUX21X1 U1262 ( .IN1(N251), .IN2(N248), .S(N308), .Q(n1140) );
  MUX41X1 U1263 ( .IN1(N254), .IN3(n776), .IN2(N242), .IN4(n777), .S0(N490), 
        .S1(N316), .Q(n864) );
  OR4X1 U1264 ( .IN1(n1063), .IN2(n1141), .IN3(n868), .IN4(n859), .Q(n1135) );
  MUX21X1 U1265 ( .IN1(n776), .IN2(n777), .S(N302), .Q(n859) );
  MUX21X1 U1266 ( .IN1(n776), .IN2(n777), .S(N361), .Q(n868) );
  INVX0 U1267 ( .INP(N248), .ZN(n777) );
  INVX0 U1268 ( .INP(N251), .ZN(n776) );
  XNOR2X1 U1269 ( .IN1(n1082), .IN2(keyinput14), .Q(n1141) );
  MUX41X1 U1270 ( .IN1(N597), .IN3(N598), .IN2(n1133), .IN4(n1134), .S0(N351), 
        .S1(n870), .Q(n1082) );
  INVX0 U1271 ( .INP(N534), .ZN(n870) );
  INVX0 U1272 ( .INP(N596), .ZN(n1133) );
  MUX21X1 U1273 ( .IN1(n1134), .IN2(N598), .S(N514), .Q(n1063) );
  INVX0 U1274 ( .INP(N595), .ZN(n1134) );
  XNOR3X1 U1275 ( .IN1(n1142), .IN2(n1143), .IN3(n1144), .Q(N7476) );
  XNOR2X1 U1276 ( .IN1(keyinput24), .IN2(n1145), .Q(n1144) );
  OA21X1 U1277 ( .IN1(n1093), .IN2(n1094), .IN3(n1146), .Q(n1145) );
  XOR2X1 U1278 ( .IN1(n1147), .IN2(keyinput16), .Q(n1146) );
  NAND2X0 U1279 ( .IN1(n1093), .IN2(n1094), .QN(n1147) );
  AO21X1 U1280 ( .IN1(N225), .IN2(N335), .IN3(n1148), .Q(n1094) );
  XOR2X1 U1281 ( .IN1(n1149), .IN2(keyinput9), .Q(n1148) );
  NAND2X0 U1282 ( .IN1(N218), .IN2(n1150), .QN(n1149) );
  INVX0 U1283 ( .INP(n1119), .ZN(n1093) );
  MUX21X1 U1284 ( .IN1(N217), .IN2(N210), .S(n1150), .Q(n1119) );
  XOR3X1 U1285 ( .IN1(n1097), .IN2(n1098), .IN3(n1151), .Q(n1143) );
  XOR2X1 U1286 ( .IN1(n1099), .IN2(n717), .Q(n1151) );
  MUX21X1 U1287 ( .IN1(N288), .IN2(N281), .S(n1150), .Q(n717) );
  MUX21X1 U1288 ( .IN1(N280), .IN2(N273), .S(n1150), .Q(n1099) );
  MUX21X1 U1289 ( .IN1(N272), .IN2(N265), .S(n1150), .Q(n1098) );
  MUX21X1 U1290 ( .IN1(N264), .IN2(N257), .S(n1150), .Q(n1097) );
  XNOR3X1 U1291 ( .IN1(n1095), .IN2(n1130), .IN3(n1152), .Q(n1142) );
  MUX21X1 U1292 ( .IN1(n1153), .IN2(n1154), .S(n1150), .Q(n1152) );
  XNOR2X1 U1293 ( .IN1(N289), .IN2(n1128), .Q(n1154) );
  XNOR2X1 U1294 ( .IN1(N292), .IN2(n1128), .Q(n1153) );
  INVX0 U1295 ( .INP(n1155), .ZN(n1128) );
  MUX21X1 U1296 ( .IN1(N209), .IN2(N206), .S(n1150), .Q(n1155) );
  MUX21X1 U1297 ( .IN1(N233), .IN2(N226), .S(n1150), .Q(n1130) );
  MUX21X1 U1298 ( .IN1(N241), .IN2(N234), .S(n1150), .Q(n1095) );
  INVX0 U1299 ( .INP(N335), .ZN(n1150) );
  OA21X1 U1300 ( .IN1(N2623), .IN2(n1156), .IN3(N141), .Q(N4740) );
  MUX21X1 U1301 ( .IN1(N82), .IN2(N80), .S(N588), .Q(n1156) );
  OA21X1 U1302 ( .IN1(N2623), .IN2(n1157), .IN3(N141), .Q(N4739) );
  MUX21X1 U1303 ( .IN1(N79), .IN2(N23), .S(N588), .Q(n1157) );
  OA21X1 U1304 ( .IN1(N2623), .IN2(n1158), .IN3(N141), .Q(N4738) );
  MUX21X1 U1305 ( .IN1(N26), .IN2(N81), .S(N588), .Q(n1158) );
  OA21X1 U1306 ( .IN1(N2623), .IN2(n1159), .IN3(N141), .Q(N4737) );
  MUX21X1 U1307 ( .IN1(N24), .IN2(N25), .S(N588), .Q(n1159) );
  NAND2X0 U1308 ( .IN1(N83), .IN2(n1160), .QN(N4279) );
  NAND2X0 U1309 ( .IN1(n1161), .IN2(n1160), .QN(N4278) );
  MUX21X1 U1310 ( .IN1(N88), .IN2(N34), .S(N588), .Q(n1161) );
  NAND2X0 U1311 ( .IN1(n1162), .IN2(n1160), .QN(N4272) );
  MUX21X1 U1312 ( .IN1(N86), .IN2(N87), .S(N588), .Q(n1162) );
  INVX0 U1313 ( .INP(N299), .ZN(N3613) );
  NAND2X0 U1314 ( .IN1(N140), .IN2(n1160), .QN(N2590) );
  INVX0 U1315 ( .INP(N2623), .ZN(n1160) );
  NAND2X0 U1316 ( .IN1(N31), .IN2(N27), .QN(N2623) );
  NAND2X0 U1317 ( .IN1(N556), .IN2(N386), .QN(N2061) );
  NAND2X0 U1318 ( .IN1(n1163), .IN2(N27), .QN(N2060) );
  INVX0 U1319 ( .INP(N591), .ZN(n1163) );
  NOR2X0 U1320 ( .IN1(N592), .IN2(n1164), .QN(N2054) );
  INVX0 U1321 ( .INP(N136), .ZN(n1164) );
  AND2X1 U1322 ( .IN1(N373), .IN2(N1), .Q(N1972) );
  INVX0 U1323 ( .INP(N559), .ZN(N1155) );
  INVX0 U1324 ( .INP(N245), .ZN(N1152) );
  AND2X1 U1325 ( .IN1(N145), .IN2(N141), .Q(N1147) );
  INVX0 U1326 ( .INP(N358), .ZN(N1145) );
  INVX0 U1327 ( .INP(N338), .ZN(N1144) );
  INVX0 U1328 ( .INP(N549), .ZN(N1141) );
  NOR2X0 U1329 ( .IN1(N1153), .IN2(N1154), .QN(N1140) );
  INVX0 U1330 ( .INP(N562), .ZN(N1154) );
  INVX0 U1331 ( .INP(N552), .ZN(N1153) );
  INVX0 U1332 ( .INP(N366), .ZN(N1139) );
  XOR2X1 U1333 ( .IN1(keyinput0), .IN2(N348), .Q(N1138) );
  INVX0 U1334 ( .INP(N545), .ZN(N1137) );
endmodule

