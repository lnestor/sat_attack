
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457;

  XNOR2X1 U289 ( .IN1(G32), .IN2(n257), .Q(G1355) );
  NOR2X0 U290 ( .IN1(n258), .IN2(n259), .QN(n257) );
  XNOR2X1 U291 ( .IN1(G31), .IN2(n260), .Q(G1354) );
  NOR2X0 U292 ( .IN1(n261), .IN2(n259), .QN(n260) );
  XNOR2X1 U293 ( .IN1(G30), .IN2(n262), .Q(G1353) );
  NOR2X0 U294 ( .IN1(n263), .IN2(n259), .QN(n262) );
  XNOR2X1 U295 ( .IN1(G29), .IN2(n264), .Q(G1352) );
  NOR2X0 U296 ( .IN1(n265), .IN2(n259), .QN(n264) );
  NAND3X0 U297 ( .IN1(n266), .IN2(n267), .IN3(n268), .QN(n259) );
  XNOR2X1 U298 ( .IN1(G28), .IN2(n269), .Q(G1351) );
  NOR2X0 U299 ( .IN1(n258), .IN2(n270), .QN(n269) );
  XNOR2X1 U300 ( .IN1(G27), .IN2(n271), .Q(G1350) );
  NOR2X0 U301 ( .IN1(n261), .IN2(n270), .QN(n271) );
  XNOR2X1 U302 ( .IN1(G26), .IN2(n272), .Q(G1349) );
  NOR2X0 U303 ( .IN1(n263), .IN2(n270), .QN(n272) );
  XNOR2X1 U304 ( .IN1(G25), .IN2(n273), .Q(G1348) );
  NOR2X0 U305 ( .IN1(n265), .IN2(n270), .QN(n273) );
  NAND4X0 U306 ( .IN1(n274), .IN2(n266), .IN3(n275), .IN4(n276), .QN(n270) );
  AND2X1 U307 ( .IN1(n277), .IN2(n267), .Q(n275) );
  XNOR2X1 U308 ( .IN1(G24), .IN2(n278), .Q(G1347) );
  NOR2X0 U309 ( .IN1(n258), .IN2(n279), .QN(n278) );
  XNOR2X1 U310 ( .IN1(G23), .IN2(n280), .Q(G1346) );
  NOR2X0 U311 ( .IN1(n261), .IN2(n279), .QN(n280) );
  XNOR2X1 U312 ( .IN1(G22), .IN2(n281), .Q(G1345) );
  NOR2X0 U313 ( .IN1(n263), .IN2(n279), .QN(n281) );
  XNOR2X1 U314 ( .IN1(G21), .IN2(n282), .Q(G1344) );
  NOR2X0 U315 ( .IN1(n265), .IN2(n279), .QN(n282) );
  NAND3X0 U316 ( .IN1(n283), .IN2(n268), .IN3(n284), .QN(n279) );
  AND3X1 U317 ( .IN1(n285), .IN2(n277), .IN3(n286), .Q(n268) );
  XNOR2X1 U318 ( .IN1(G20), .IN2(n287), .Q(G1343) );
  NOR2X0 U319 ( .IN1(n258), .IN2(n288), .QN(n287) );
  XNOR2X1 U320 ( .IN1(G19), .IN2(n289), .Q(G1342) );
  NOR2X0 U321 ( .IN1(n261), .IN2(n288), .QN(n289) );
  XNOR2X1 U322 ( .IN1(G18), .IN2(n290), .Q(G1341) );
  NOR2X0 U323 ( .IN1(n263), .IN2(n288), .QN(n290) );
  XNOR2X1 U324 ( .IN1(G17), .IN2(n291), .Q(G1340) );
  NOR2X0 U325 ( .IN1(n265), .IN2(n288), .QN(n291) );
  NAND4X0 U326 ( .IN1(n283), .IN2(n292), .IN3(n276), .IN4(n277), .QN(n288) );
  NAND2X0 U327 ( .IN1(n293), .IN2(n294), .QN(n277) );
  OR3X1 U328 ( .IN1(n295), .IN2(n296), .IN3(n297), .Q(n294) );
  OR3X1 U329 ( .IN1(n298), .IN2(n299), .IN3(n300), .Q(n293) );
  XNOR2X1 U330 ( .IN1(G16), .IN2(n301), .Q(G1339) );
  NOR2X0 U331 ( .IN1(n302), .IN2(n276), .QN(n301) );
  XNOR2X1 U332 ( .IN1(G15), .IN2(n303), .Q(G1338) );
  NOR2X0 U333 ( .IN1(n302), .IN2(n285), .QN(n303) );
  XNOR2X1 U334 ( .IN1(G14), .IN2(n304), .Q(G1337) );
  NOR2X0 U335 ( .IN1(n283), .IN2(n302), .QN(n304) );
  XOR2X1 U336 ( .IN1(n305), .IN2(G12), .Q(G1335) );
  NAND2X0 U337 ( .IN1(n306), .IN2(n286), .QN(n305) );
  XOR2X1 U338 ( .IN1(n307), .IN2(G11), .Q(G1334) );
  NAND2X0 U339 ( .IN1(n306), .IN2(n274), .QN(n307) );
  XOR2X1 U340 ( .IN1(n308), .IN2(G10), .Q(G1333) );
  NAND2X0 U341 ( .IN1(n306), .IN2(n266), .QN(n308) );
  XOR2X1 U342 ( .IN1(n309), .IN2(G9), .Q(G1332) );
  NAND2X0 U343 ( .IN1(n306), .IN2(n284), .QN(n309) );
  AND4X1 U344 ( .IN1(n295), .IN2(n310), .IN3(n298), .IN4(n258), .Q(n306) );
  XNOR2X1 U345 ( .IN1(G8), .IN2(n311), .Q(G1331) );
  NOR2X0 U346 ( .IN1(n276), .IN2(n312), .QN(n311) );
  XNOR2X1 U347 ( .IN1(G7), .IN2(n313), .Q(G1330) );
  NOR2X0 U348 ( .IN1(n285), .IN2(n312), .QN(n313) );
  XNOR2X1 U349 ( .IN1(G6), .IN2(n314), .Q(G1329) );
  NOR2X0 U350 ( .IN1(n283), .IN2(n312), .QN(n314) );
  XNOR2X1 U351 ( .IN1(G5), .IN2(n315), .Q(G1328) );
  NOR2X0 U352 ( .IN1(n267), .IN2(n312), .QN(n315) );
  NAND4X0 U353 ( .IN1(n297), .IN2(n316), .IN3(n317), .IN4(n300), .QN(n312) );
  NOR2X0 U354 ( .IN1(n298), .IN2(n295), .QN(n317) );
  XNOR2X1 U355 ( .IN1(G4), .IN2(n318), .Q(G1327) );
  NOR2X0 U356 ( .IN1(n276), .IN2(n319), .QN(n318) );
  INVX0 U357 ( .INP(n286), .ZN(n276) );
  XNOR2X1 U358 ( .IN1(G3), .IN2(n320), .Q(G1326) );
  NOR2X0 U359 ( .IN1(n285), .IN2(n319), .QN(n320) );
  XNOR2X1 U360 ( .IN1(G2), .IN2(n321), .Q(G1325) );
  NOR2X0 U361 ( .IN1(n283), .IN2(n319), .QN(n321) );
  XNOR2X1 U362 ( .IN1(G1), .IN2(n322), .Q(G1324) );
  NOR2X0 U363 ( .IN1(n267), .IN2(n319), .QN(n322) );
  NAND4X0 U364 ( .IN1(n316), .IN2(n296), .IN3(n258), .IN4(n263), .QN(n319) );
  NOR2X0 U365 ( .IN1(n261), .IN2(n265), .QN(n296) );
  XOR3X1 U366 ( .IN1(keyinput31), .IN2(keyinput30), .IN3(n323), .Q(G1336) );
  NOR2X0 U367 ( .IN1(n324), .IN2(n325), .QN(n323) );
  XOR2X1 U368 ( .IN1(keyinput28), .IN2(n326), .Q(n325) );
  NOR2X0 U369 ( .IN1(n327), .IN2(n328), .QN(n326) );
  XOR2X1 U370 ( .IN1(keyinput29), .IN2(n329), .Q(n324) );
  NOR2X0 U371 ( .IN1(n327), .IN2(n330), .QN(n329) );
  XOR2X1 U372 ( .IN1(n331), .IN2(keyinput27), .Q(n327) );
  OR2X1 U373 ( .IN1(n330), .IN2(n328), .Q(n331) );
  XNOR2X1 U374 ( .IN1(n332), .IN2(keyinput26), .Q(n330) );
  OR2X1 U375 ( .IN1(n267), .IN2(n302), .Q(n332) );
  XOR2X1 U376 ( .IN1(n333), .IN2(keyinput25), .Q(n302) );
  NAND3X0 U377 ( .IN1(n310), .IN2(n261), .IN3(n299), .QN(n333) );
  NOR2X0 U378 ( .IN1(n263), .IN2(n258), .QN(n299) );
  INVX0 U379 ( .INP(n297), .ZN(n258) );
  MUX21X1 U380 ( .IN1(n334), .IN2(n335), .S(n336), .Q(n297) );
  XOR3X1 U381 ( .IN1(G24), .IN2(G20), .IN3(n337), .Q(n336) );
  XOR2X1 U382 ( .IN1(G32), .IN2(G28), .Q(n337) );
  NAND2X0 U383 ( .IN1(n338), .IN2(n339), .QN(n335) );
  AND2X1 U384 ( .IN1(n339), .IN2(n338), .Q(n334) );
  NAND3X0 U385 ( .IN1(G41), .IN2(n340), .IN3(G40), .QN(n338) );
  AO21X1 U386 ( .IN1(G40), .IN2(G41), .IN3(n340), .Q(n339) );
  XOR2X1 U387 ( .IN1(n341), .IN2(n342), .Q(n340) );
  INVX0 U388 ( .INP(n295), .ZN(n263) );
  MUX21X1 U389 ( .IN1(n343), .IN2(n344), .S(n345), .Q(n295) );
  XNOR3X1 U390 ( .IN1(n346), .IN2(G18), .IN3(n347), .Q(n345) );
  XNOR2X1 U391 ( .IN1(n348), .IN2(G26), .Q(n347) );
  INVX0 U392 ( .INP(G22), .ZN(n346) );
  NAND2X0 U393 ( .IN1(n349), .IN2(n350), .QN(n344) );
  AND2X1 U394 ( .IN1(n350), .IN2(n349), .Q(n343) );
  NAND3X0 U395 ( .IN1(G41), .IN2(n351), .IN3(G38), .QN(n349) );
  AO21X1 U396 ( .IN1(G38), .IN2(G41), .IN3(n351), .Q(n350) );
  XOR2X1 U397 ( .IN1(n341), .IN2(n352), .Q(n351) );
  XNOR3X1 U398 ( .IN1(G14), .IN2(G13), .IN3(n353), .Q(n341) );
  XNOR3X1 U399 ( .IN1(keyinput4), .IN2(G16), .IN3(G15), .Q(n353) );
  INVX0 U400 ( .INP(n298), .ZN(n261) );
  MUX21X1 U401 ( .IN1(n354), .IN2(n355), .S(n356), .Q(n298) );
  XNOR3X1 U402 ( .IN1(n357), .IN2(G19), .IN3(n358), .Q(n356) );
  OA21X1 U403 ( .IN1(G27), .IN2(G31), .IN3(n359), .Q(n358) );
  XOR2X1 U404 ( .IN1(keyinput1), .IN2(n360), .Q(n359) );
  AND2X1 U405 ( .IN1(G27), .IN2(G31), .Q(n360) );
  INVX0 U406 ( .INP(G23), .ZN(n357) );
  NAND2X0 U407 ( .IN1(n361), .IN2(n362), .QN(n355) );
  AND2X1 U408 ( .IN1(n362), .IN2(n361), .Q(n354) );
  NAND3X0 U409 ( .IN1(G39), .IN2(n363), .IN3(G41), .QN(n361) );
  AO21X1 U410 ( .IN1(G41), .IN2(G39), .IN3(n363), .Q(n362) );
  XOR2X1 U411 ( .IN1(n364), .IN2(n352), .Q(n363) );
  XNOR3X1 U412 ( .IN1(G11), .IN2(G10), .IN3(n365), .Q(n352) );
  XNOR2X1 U413 ( .IN1(G12), .IN2(G9), .Q(n365) );
  AND2X1 U414 ( .IN1(n316), .IN2(n265), .Q(n310) );
  INVX0 U415 ( .INP(n300), .ZN(n265) );
  MUX21X1 U416 ( .IN1(n366), .IN2(n367), .S(n368), .Q(n300) );
  XOR3X1 U417 ( .IN1(G21), .IN2(G17), .IN3(n369), .Q(n368) );
  XNOR2X1 U418 ( .IN1(n370), .IN2(G25), .Q(n369) );
  NAND2X0 U419 ( .IN1(n371), .IN2(n372), .QN(n367) );
  AND2X1 U420 ( .IN1(n372), .IN2(n371), .Q(n366) );
  NAND3X0 U421 ( .IN1(G41), .IN2(n373), .IN3(G37), .QN(n371) );
  AO21X1 U422 ( .IN1(G37), .IN2(G41), .IN3(n373), .Q(n372) );
  XOR2X1 U423 ( .IN1(n342), .IN2(n364), .Q(n373) );
  XNOR3X1 U424 ( .IN1(G2), .IN2(G1), .IN3(n374), .Q(n364) );
  XNOR2X1 U425 ( .IN1(G3), .IN2(G4), .Q(n374) );
  XNOR3X1 U426 ( .IN1(G6), .IN2(G5), .IN3(n375), .Q(n342) );
  XNOR2X1 U427 ( .IN1(G7), .IN2(G8), .Q(n375) );
  XOR2X1 U428 ( .IN1(n376), .IN2(keyinput24), .Q(n316) );
  AO222X1 U429 ( .IN1(n377), .IN2(n285), .IN3(n378), .IN4(n283), .IN5(
        keyinput23), .IN6(n379), .Q(n376) );
  NAND3X0 U430 ( .IN1(n285), .IN2(n267), .IN3(n380), .QN(n379) );
  XNOR2X1 U431 ( .IN1(keyinput22), .IN2(n283), .Q(n380) );
  INVX0 U432 ( .INP(n266), .ZN(n283) );
  NOR2X0 U433 ( .IN1(n292), .IN2(n286), .QN(n378) );
  NOR2X0 U434 ( .IN1(n267), .IN2(n285), .QN(n292) );
  INVX0 U435 ( .INP(n274), .ZN(n285) );
  MUX21X1 U436 ( .IN1(n381), .IN2(n382), .S(n383), .Q(n274) );
  XNOR3X1 U437 ( .IN1(n384), .IN2(G11), .IN3(n385), .Q(n383) );
  XNOR2X1 U438 ( .IN1(n386), .IN2(G3), .Q(n385) );
  INVX0 U439 ( .INP(G7), .ZN(n386) );
  INVX0 U440 ( .INP(G15), .ZN(n384) );
  NAND2X0 U441 ( .IN1(n387), .IN2(n388), .QN(n382) );
  AND2X1 U442 ( .IN1(n388), .IN2(n387), .Q(n381) );
  NAND3X0 U443 ( .IN1(G41), .IN2(n389), .IN3(G35), .QN(n387) );
  AO21X1 U444 ( .IN1(G35), .IN2(G41), .IN3(n389), .Q(n388) );
  XOR2X1 U445 ( .IN1(n390), .IN2(n391), .Q(n389) );
  NOR2X0 U446 ( .IN1(n392), .IN2(n284), .QN(n377) );
  OA21X1 U447 ( .IN1(keyinput23), .IN2(n393), .IN3(n286), .Q(n392) );
  MUX21X1 U448 ( .IN1(n394), .IN2(n395), .S(n396), .Q(n286) );
  XOR3X1 U449 ( .IN1(G16), .IN2(G12), .IN3(n397), .Q(n396) );
  XOR2X1 U450 ( .IN1(G8), .IN2(G4), .Q(n397) );
  NAND2X0 U451 ( .IN1(n398), .IN2(n399), .QN(n395) );
  AND2X1 U452 ( .IN1(n399), .IN2(n398), .Q(n394) );
  NAND3X0 U453 ( .IN1(G41), .IN2(n400), .IN3(G36), .QN(n398) );
  AO21X1 U454 ( .IN1(G36), .IN2(G41), .IN3(n400), .Q(n399) );
  XOR2X1 U455 ( .IN1(n401), .IN2(n402), .Q(n400) );
  XNOR2X1 U456 ( .IN1(n266), .IN2(keyinput22), .Q(n393) );
  XNOR2X1 U457 ( .IN1(n403), .IN2(keyinput21), .Q(n266) );
  NAND2X0 U458 ( .IN1(n404), .IN2(n405), .QN(n403) );
  XOR2X1 U459 ( .IN1(keyinput19), .IN2(n406), .Q(n405) );
  NOR2X0 U460 ( .IN1(n407), .IN2(n408), .QN(n406) );
  XOR2X1 U461 ( .IN1(keyinput18), .IN2(n409), .Q(n408) );
  XOR2X1 U462 ( .IN1(n410), .IN2(keyinput20), .Q(n404) );
  NAND2X0 U463 ( .IN1(n411), .IN2(n412), .QN(n410) );
  INVX0 U464 ( .INP(n413), .ZN(n412) );
  XNOR2X1 U465 ( .IN1(keyinput18), .IN2(n409), .Q(n411) );
  NOR2X0 U466 ( .IN1(n413), .IN2(n407), .QN(n409) );
  XNOR3X1 U467 ( .IN1(n414), .IN2(G10), .IN3(n415), .Q(n407) );
  XNOR2X1 U468 ( .IN1(G2), .IN2(G6), .Q(n415) );
  INVX0 U469 ( .INP(G14), .ZN(n414) );
  XNOR2X1 U470 ( .IN1(n416), .IN2(keyinput17), .Q(n413) );
  NAND2X0 U471 ( .IN1(n417), .IN2(n418), .QN(n416) );
  XNOR2X1 U472 ( .IN1(n419), .IN2(keyinput15), .Q(n418) );
  NAND3X0 U473 ( .IN1(G41), .IN2(n420), .IN3(G34), .QN(n419) );
  XOR2X1 U474 ( .IN1(n421), .IN2(keyinput16), .Q(n417) );
  NAND2X0 U475 ( .IN1(n420), .IN2(n422), .QN(n421) );
  XNOR2X1 U476 ( .IN1(n423), .IN2(keyinput14), .Q(n420) );
  NAND3X0 U477 ( .IN1(G41), .IN2(n422), .IN3(G34), .QN(n423) );
  XNOR2X1 U478 ( .IN1(n424), .IN2(keyinput13), .Q(n422) );
  NAND2X0 U479 ( .IN1(n425), .IN2(n426), .QN(n424) );
  XOR2X1 U480 ( .IN1(keyinput12), .IN2(n427), .Q(n426) );
  AND2X1 U481 ( .IN1(n402), .IN2(n428), .Q(n427) );
  XOR2X1 U482 ( .IN1(n429), .IN2(keyinput11), .Q(n425) );
  NAND2X0 U483 ( .IN1(n428), .IN2(n391), .QN(n429) );
  XOR2X1 U484 ( .IN1(n430), .IN2(keyinput10), .Q(n428) );
  NAND2X0 U485 ( .IN1(n391), .IN2(n402), .QN(n430) );
  XNOR2X1 U486 ( .IN1(n431), .IN2(keyinput9), .Q(n402) );
  NAND2X0 U487 ( .IN1(n432), .IN2(n433), .QN(n431) );
  XOR2X1 U488 ( .IN1(n434), .IN2(keyinput8), .Q(n433) );
  NAND2X0 U489 ( .IN1(n435), .IN2(n436), .QN(n434) );
  XOR2X1 U490 ( .IN1(n437), .IN2(keyinput7), .Q(n432) );
  NAND2X0 U491 ( .IN1(n438), .IN2(n435), .QN(n437) );
  XNOR2X1 U492 ( .IN1(n439), .IN2(keyinput6), .Q(n435) );
  NAND2X0 U493 ( .IN1(n438), .IN2(n436), .QN(n439) );
  XOR2X1 U494 ( .IN1(G32), .IN2(G31), .Q(n436) );
  XOR2X1 U495 ( .IN1(n440), .IN2(keyinput5), .Q(n438) );
  NAND2X0 U496 ( .IN1(n441), .IN2(n442), .QN(n440) );
  XOR2X1 U497 ( .IN1(keyinput2), .IN2(n443), .Q(n442) );
  NOR2X0 U498 ( .IN1(n370), .IN2(n444), .QN(n443) );
  INVX0 U499 ( .INP(G29), .ZN(n370) );
  XOR2X1 U500 ( .IN1(n445), .IN2(keyinput3), .Q(n441) );
  OR2X1 U501 ( .IN1(n444), .IN2(n348), .Q(n445) );
  INVX0 U502 ( .INP(G30), .ZN(n348) );
  XNOR2X1 U503 ( .IN1(n446), .IN2(keyinput0), .Q(n444) );
  NAND2X0 U504 ( .IN1(G30), .IN2(G29), .QN(n446) );
  XNOR3X1 U505 ( .IN1(G26), .IN2(G25), .IN3(n447), .Q(n391) );
  XNOR2X1 U506 ( .IN1(G28), .IN2(G27), .Q(n447) );
  INVX0 U507 ( .INP(n284), .ZN(n267) );
  MUX21X1 U508 ( .IN1(n448), .IN2(n449), .S(n450), .Q(n284) );
  XNOR3X1 U509 ( .IN1(n328), .IN2(G1), .IN3(n451), .Q(n450) );
  XNOR2X1 U510 ( .IN1(G9), .IN2(n452), .Q(n451) );
  INVX0 U511 ( .INP(G5), .ZN(n452) );
  INVX0 U512 ( .INP(G13), .ZN(n328) );
  NAND2X0 U513 ( .IN1(n453), .IN2(n454), .QN(n449) );
  AND2X1 U514 ( .IN1(n454), .IN2(n453), .Q(n448) );
  NAND3X0 U515 ( .IN1(G41), .IN2(n455), .IN3(G33), .QN(n453) );
  AO21X1 U516 ( .IN1(G33), .IN2(G41), .IN3(n455), .Q(n454) );
  XOR2X1 U517 ( .IN1(n390), .IN2(n401), .Q(n455) );
  XNOR3X1 U518 ( .IN1(G22), .IN2(G21), .IN3(n456), .Q(n401) );
  XNOR2X1 U519 ( .IN1(G23), .IN2(G24), .Q(n456) );
  XNOR3X1 U520 ( .IN1(G18), .IN2(G17), .IN3(n457), .Q(n390) );
  XNOR2X1 U521 ( .IN1(G19), .IN2(G20), .Q(n457) );
endmodule

