
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168;

  XOR3X1 U613 ( .IN1(keyinput253), .IN2(keyinput235), .IN3(n590), .Q(G1343) );
  NOR2X0 U614 ( .IN1(n591), .IN2(n592), .QN(n590) );
  XOR2X1 U615 ( .IN1(keyinput213), .IN2(n593), .Q(n592) );
  AND2X1 U616 ( .IN1(G20), .IN2(n594), .Q(n593) );
  XOR2X1 U617 ( .IN1(n595), .IN2(keyinput214), .Q(n591) );
  NAND2X0 U618 ( .IN1(n594), .IN2(n596), .QN(n595) );
  XOR2X1 U619 ( .IN1(n597), .IN2(keyinput180), .Q(n594) );
  NAND2X0 U620 ( .IN1(G20), .IN2(n596), .QN(n597) );
  XNOR2X1 U621 ( .IN1(n598), .IN2(keyinput161), .Q(n596) );
  NAND2X0 U622 ( .IN1(n599), .IN2(n600), .QN(n598) );
  XOR3X1 U623 ( .IN1(keyinput252), .IN2(keyinput234), .IN3(n601), .Q(G1342) );
  NAND2X0 U624 ( .IN1(n602), .IN2(n603), .QN(n601) );
  XOR2X1 U625 ( .IN1(keyinput211), .IN2(n604), .Q(n603) );
  NOR2X0 U626 ( .IN1(n605), .IN2(n606), .QN(n604) );
  XOR2X1 U627 ( .IN1(keyinput212), .IN2(n607), .Q(n602) );
  NOR2X0 U628 ( .IN1(n608), .IN2(n606), .QN(n607) );
  XNOR2X1 U629 ( .IN1(n609), .IN2(keyinput179), .Q(n606) );
  OR2X1 U630 ( .IN1(n608), .IN2(n605), .Q(n609) );
  INVX0 U631 ( .INP(G19), .ZN(n605) );
  XNOR2X1 U632 ( .IN1(n610), .IN2(keyinput160), .Q(n608) );
  NAND2X0 U633 ( .IN1(n611), .IN2(n599), .QN(n610) );
  XOR3X1 U634 ( .IN1(keyinput249), .IN2(keyinput231), .IN3(n612), .Q(G1339) );
  NOR2X0 U635 ( .IN1(n613), .IN2(n614), .QN(n612) );
  XOR2X1 U636 ( .IN1(keyinput205), .IN2(n615), .Q(n614) );
  NOR2X0 U637 ( .IN1(n616), .IN2(n617), .QN(n615) );
  XOR2X1 U638 ( .IN1(keyinput206), .IN2(n618), .Q(n613) );
  NOR2X0 U639 ( .IN1(n619), .IN2(n616), .QN(n618) );
  XOR2X1 U640 ( .IN1(n620), .IN2(keyinput176), .Q(n616) );
  OR2X1 U641 ( .IN1(n617), .IN2(n619), .Q(n620) );
  XOR2X1 U642 ( .IN1(n621), .IN2(keyinput157), .Q(n619) );
  NAND2X0 U643 ( .IN1(n622), .IN2(n623), .QN(n621) );
  XOR3X1 U644 ( .IN1(keyinput244), .IN2(keyinput226), .IN3(n624), .Q(G1334) );
  NAND2X0 U645 ( .IN1(n625), .IN2(n626), .QN(n624) );
  XOR2X1 U646 ( .IN1(keyinput195), .IN2(n627), .Q(n626) );
  NOR2X0 U647 ( .IN1(n628), .IN2(n629), .QN(n627) );
  XOR2X1 U648 ( .IN1(keyinput196), .IN2(n630), .Q(n625) );
  NOR2X0 U649 ( .IN1(n628), .IN2(n631), .QN(n630) );
  XOR2X1 U650 ( .IN1(n632), .IN2(keyinput171), .Q(n628) );
  OR2X1 U651 ( .IN1(n631), .IN2(n629), .Q(n632) );
  INVX0 U652 ( .INP(G11), .ZN(n629) );
  XNOR2X1 U653 ( .IN1(n633), .IN2(keyinput152), .Q(n631) );
  NAND2X0 U654 ( .IN1(n634), .IN2(n635), .QN(n633) );
  XOR3X1 U655 ( .IN1(keyinput241), .IN2(keyinput223), .IN3(n636), .Q(G1327) );
  NAND2X0 U656 ( .IN1(n637), .IN2(n638), .QN(n636) );
  XOR2X1 U657 ( .IN1(n639), .IN2(keyinput189), .Q(n638) );
  NAND2X0 U658 ( .IN1(n640), .IN2(G4), .QN(n639) );
  XOR2X1 U659 ( .IN1(n641), .IN2(keyinput190), .Q(n637) );
  NAND2X0 U660 ( .IN1(n640), .IN2(n642), .QN(n641) );
  XOR2X1 U661 ( .IN1(n643), .IN2(keyinput168), .Q(n640) );
  NAND2X0 U662 ( .IN1(n642), .IN2(G4), .QN(n643) );
  XOR2X1 U663 ( .IN1(n644), .IN2(keyinput149), .Q(n642) );
  NAND2X0 U664 ( .IN1(n645), .IN2(n623), .QN(n644) );
  XOR3X1 U665 ( .IN1(keyinput240), .IN2(keyinput222), .IN3(n646), .Q(G1326) );
  NAND2X0 U666 ( .IN1(n647), .IN2(n648), .QN(n646) );
  XOR2X1 U667 ( .IN1(keyinput188), .IN2(n649), .Q(n648) );
  AND2X1 U668 ( .IN1(n650), .IN2(n651), .Q(n649) );
  XOR2X1 U669 ( .IN1(n652), .IN2(keyinput187), .Q(n647) );
  NAND2X0 U670 ( .IN1(n651), .IN2(G3), .QN(n652) );
  XOR2X1 U671 ( .IN1(n653), .IN2(keyinput167), .Q(n651) );
  NAND2X0 U672 ( .IN1(G3), .IN2(n650), .QN(n653) );
  XNOR2X1 U673 ( .IN1(n654), .IN2(keyinput148), .Q(n650) );
  NAND2X0 U674 ( .IN1(n645), .IN2(n635), .QN(n654) );
  XOR3X1 U675 ( .IN1(keyinput238), .IN2(keyinput220), .IN3(n655), .Q(G1324) );
  NOR2X0 U676 ( .IN1(n656), .IN2(n657), .QN(n655) );
  XOR2X1 U677 ( .IN1(n658), .IN2(keyinput184), .Q(n657) );
  NAND2X0 U678 ( .IN1(n659), .IN2(n660), .QN(n658) );
  XOR2X1 U679 ( .IN1(n661), .IN2(keyinput183), .Q(n656) );
  NAND2X0 U680 ( .IN1(G1), .IN2(n659), .QN(n661) );
  XNOR2X1 U681 ( .IN1(n662), .IN2(keyinput165), .Q(n659) );
  NAND2X0 U682 ( .IN1(G1), .IN2(n660), .QN(n662) );
  XNOR2X1 U683 ( .IN1(n663), .IN2(keyinput146), .Q(n660) );
  NAND2X0 U684 ( .IN1(n645), .IN2(n664), .QN(n663) );
  XOR3X1 U685 ( .IN1(keyinput164), .IN2(G32), .IN3(n665), .Q(G1355) );
  NOR2X0 U686 ( .IN1(n666), .IN2(n667), .QN(n665) );
  NOR2X0 U687 ( .IN1(n668), .IN2(n669), .QN(G1354) );
  XOR2X1 U688 ( .IN1(n670), .IN2(keyinput219), .Q(n669) );
  NAND3X0 U689 ( .IN1(n611), .IN2(n671), .IN3(n672), .QN(n670) );
  OA21X1 U690 ( .IN1(n673), .IN2(n667), .IN3(G31), .Q(n668) );
  XOR2X1 U691 ( .IN1(n674), .IN2(G30), .Q(G1353) );
  NAND2X0 U692 ( .IN1(n672), .IN2(n675), .QN(n674) );
  XOR2X1 U693 ( .IN1(n676), .IN2(G29), .Q(G1352) );
  NAND2X0 U694 ( .IN1(n672), .IN2(n677), .QN(n676) );
  INVX0 U695 ( .INP(n667), .ZN(n672) );
  NAND4X0 U696 ( .IN1(n623), .IN2(n678), .IN3(n679), .IN4(n680), .QN(n667) );
  NOR2X0 U697 ( .IN1(n681), .IN2(n664), .QN(n679) );
  XNOR2X1 U698 ( .IN1(G28), .IN2(n682), .Q(G1351) );
  NOR2X0 U699 ( .IN1(n666), .IN2(n683), .QN(n682) );
  XNOR2X1 U700 ( .IN1(G27), .IN2(n684), .Q(G1350) );
  NOR2X0 U701 ( .IN1(n673), .IN2(n683), .QN(n684) );
  XOR2X1 U702 ( .IN1(n685), .IN2(n686), .Q(G1349) );
  NOR2X0 U703 ( .IN1(n687), .IN2(n683), .QN(n686) );
  XOR2X1 U704 ( .IN1(n688), .IN2(n689), .Q(G1348) );
  NOR2X0 U705 ( .IN1(n690), .IN2(n683), .QN(n689) );
  NAND4X0 U706 ( .IN1(n680), .IN2(n691), .IN3(n635), .IN4(n692), .QN(n683) );
  XOR2X1 U707 ( .IN1(n693), .IN2(n694), .Q(G1346) );
  NOR2X0 U708 ( .IN1(n695), .IN2(n673), .QN(n694) );
  INVX0 U709 ( .INP(n611), .ZN(n673) );
  XOR2X1 U710 ( .IN1(n696), .IN2(n697), .Q(G1344) );
  NOR2X0 U711 ( .IN1(n695), .IN2(n690), .QN(n697) );
  XOR2X1 U712 ( .IN1(n698), .IN2(G8), .Q(G1331) );
  NAND2X0 U713 ( .IN1(n699), .IN2(n623), .QN(n698) );
  XOR2X1 U714 ( .IN1(n700), .IN2(G7), .Q(G1330) );
  NAND2X0 U715 ( .IN1(n699), .IN2(n635), .QN(n700) );
  XOR2X1 U716 ( .IN1(n701), .IN2(G6), .Q(G1329) );
  NAND2X0 U717 ( .IN1(n699), .IN2(n680), .QN(n701) );
  XOR2X1 U718 ( .IN1(n702), .IN2(G5), .Q(G1328) );
  NAND2X0 U719 ( .IN1(n699), .IN2(n664), .QN(n702) );
  AND2X1 U720 ( .IN1(n703), .IN2(n704), .Q(n699) );
  XOR3X1 U721 ( .IN1(keyinput255), .IN2(keyinput237), .IN3(n705), .Q(G1347) );
  NAND2X0 U722 ( .IN1(n706), .IN2(n707), .QN(n705) );
  XOR2X1 U723 ( .IN1(keyinput217), .IN2(n708), .Q(n707) );
  NOR2X0 U724 ( .IN1(n709), .IN2(n710), .QN(n708) );
  XOR2X1 U725 ( .IN1(keyinput218), .IN2(n711), .Q(n706) );
  NOR2X0 U726 ( .IN1(n712), .IN2(n709), .QN(n711) );
  XOR2X1 U727 ( .IN1(n713), .IN2(keyinput182), .Q(n709) );
  OR2X1 U728 ( .IN1(n710), .IN2(n712), .Q(n713) );
  XOR2X1 U729 ( .IN1(n714), .IN2(keyinput163), .Q(n712) );
  NAND2X0 U730 ( .IN1(n600), .IN2(n715), .QN(n714) );
  XOR3X1 U731 ( .IN1(keyinput254), .IN2(keyinput236), .IN3(n716), .Q(G1345) );
  NAND2X0 U732 ( .IN1(n717), .IN2(n718), .QN(n716) );
  XOR2X1 U733 ( .IN1(keyinput215), .IN2(n719), .Q(n718) );
  NOR2X0 U734 ( .IN1(n720), .IN2(n721), .QN(n719) );
  XOR2X1 U735 ( .IN1(keyinput216), .IN2(n722), .Q(n717) );
  NOR2X0 U736 ( .IN1(n720), .IN2(n723), .QN(n722) );
  XOR2X1 U737 ( .IN1(n724), .IN2(keyinput181), .Q(n720) );
  OR2X1 U738 ( .IN1(n723), .IN2(n721), .Q(n724) );
  XNOR2X1 U739 ( .IN1(n725), .IN2(keyinput162), .Q(n723) );
  NAND2X0 U740 ( .IN1(n675), .IN2(n715), .QN(n725) );
  INVX0 U741 ( .INP(n695), .ZN(n715) );
  XOR2X1 U742 ( .IN1(n726), .IN2(keyinput145), .Q(n695) );
  NAND4X0 U743 ( .IN1(n664), .IN2(n727), .IN3(n623), .IN4(n692), .QN(n726) );
  XOR3X1 U744 ( .IN1(keyinput251), .IN2(keyinput233), .IN3(n728), .Q(G1341) );
  NOR2X0 U745 ( .IN1(n729), .IN2(n730), .QN(n728) );
  XOR2X1 U746 ( .IN1(n731), .IN2(keyinput210), .Q(n730) );
  NAND2X0 U747 ( .IN1(n732), .IN2(n733), .QN(n731) );
  XOR2X1 U748 ( .IN1(n734), .IN2(keyinput209), .Q(n729) );
  NAND2X0 U749 ( .IN1(G18), .IN2(n733), .QN(n734) );
  XNOR2X1 U750 ( .IN1(n735), .IN2(keyinput178), .Q(n733) );
  NAND2X0 U751 ( .IN1(n732), .IN2(G18), .QN(n735) );
  XOR2X1 U752 ( .IN1(n736), .IN2(keyinput159), .Q(n732) );
  NAND2X0 U753 ( .IN1(n599), .IN2(n675), .QN(n736) );
  XOR3X1 U754 ( .IN1(keyinput250), .IN2(keyinput232), .IN3(n737), .Q(G1340) );
  NOR2X0 U755 ( .IN1(n738), .IN2(n739), .QN(n737) );
  XOR2X1 U756 ( .IN1(n740), .IN2(keyinput208), .Q(n739) );
  NAND2X0 U757 ( .IN1(n741), .IN2(n742), .QN(n740) );
  XOR2X1 U758 ( .IN1(n743), .IN2(keyinput207), .Q(n738) );
  NAND2X0 U759 ( .IN1(n741), .IN2(G17), .QN(n743) );
  XOR2X1 U760 ( .IN1(n744), .IN2(keyinput177), .Q(n741) );
  NAND2X0 U761 ( .IN1(n742), .IN2(G17), .QN(n744) );
  XOR2X1 U762 ( .IN1(n745), .IN2(keyinput158), .Q(n742) );
  NAND2X0 U763 ( .IN1(n677), .IN2(n599), .QN(n745) );
  XOR2X1 U764 ( .IN1(n746), .IN2(keyinput144), .Q(n599) );
  NAND4X0 U765 ( .IN1(n747), .IN2(n664), .IN3(n748), .IN4(n749), .QN(n746) );
  XNOR2X1 U766 ( .IN1(keyinput133), .IN2(n680), .Q(n749) );
  NOR2X0 U767 ( .IN1(n681), .IN2(n678), .QN(n748) );
  INVX0 U768 ( .INP(n692), .ZN(n681) );
  NAND2X0 U769 ( .IN1(n750), .IN2(n751), .QN(n692) );
  OAI221X1 U770 ( .IN1(n687), .IN2(n752), .IN3(n666), .IN4(n704), .IN5(n690), 
        .QN(n751) );
  XOR2X1 U771 ( .IN1(n753), .IN2(keyinput139), .Q(n750) );
  NAND2X0 U772 ( .IN1(n752), .IN2(n687), .QN(n753) );
  NOR2X0 U773 ( .IN1(n600), .IN2(n611), .QN(n752) );
  XOR2X1 U774 ( .IN1(n623), .IN2(keyinput134), .Q(n747) );
  XOR3X1 U775 ( .IN1(keyinput248), .IN2(keyinput230), .IN3(n754), .Q(G1338) );
  NOR2X0 U776 ( .IN1(n755), .IN2(n756), .QN(n754) );
  XOR2X1 U777 ( .IN1(n757), .IN2(keyinput204), .Q(n756) );
  NAND2X0 U778 ( .IN1(n758), .IN2(n759), .QN(n757) );
  XOR2X1 U779 ( .IN1(n760), .IN2(keyinput203), .Q(n755) );
  NAND2X0 U780 ( .IN1(n758), .IN2(G15), .QN(n760) );
  XOR2X1 U781 ( .IN1(n761), .IN2(keyinput175), .Q(n758) );
  NAND2X0 U782 ( .IN1(G15), .IN2(n759), .QN(n761) );
  XNOR2X1 U783 ( .IN1(n762), .IN2(keyinput156), .Q(n759) );
  NAND2X0 U784 ( .IN1(n622), .IN2(n635), .QN(n762) );
  XOR3X1 U785 ( .IN1(keyinput247), .IN2(keyinput229), .IN3(n763), .Q(G1337) );
  NOR2X0 U786 ( .IN1(n764), .IN2(n765), .QN(n763) );
  XOR2X1 U787 ( .IN1(n766), .IN2(keyinput202), .Q(n765) );
  NAND2X0 U788 ( .IN1(n767), .IN2(n768), .QN(n766) );
  XOR2X1 U789 ( .IN1(n769), .IN2(keyinput201), .Q(n764) );
  NAND2X0 U790 ( .IN1(G14), .IN2(n768), .QN(n769) );
  XNOR2X1 U791 ( .IN1(n770), .IN2(keyinput174), .Q(n768) );
  NAND2X0 U792 ( .IN1(n767), .IN2(G14), .QN(n770) );
  XOR2X1 U793 ( .IN1(n771), .IN2(keyinput155), .Q(n767) );
  NAND2X0 U794 ( .IN1(n622), .IN2(n680), .QN(n771) );
  XOR3X1 U795 ( .IN1(keyinput246), .IN2(keyinput228), .IN3(n772), .Q(G1336) );
  NOR2X0 U796 ( .IN1(n773), .IN2(n774), .QN(n772) );
  XOR2X1 U797 ( .IN1(keyinput199), .IN2(n775), .Q(n774) );
  NOR2X0 U798 ( .IN1(n776), .IN2(n777), .QN(n775) );
  XOR2X1 U799 ( .IN1(keyinput200), .IN2(n778), .Q(n773) );
  NOR2X0 U800 ( .IN1(n779), .IN2(n777), .QN(n778) );
  XNOR2X1 U801 ( .IN1(n780), .IN2(keyinput173), .Q(n777) );
  OR2X1 U802 ( .IN1(n779), .IN2(n776), .Q(n780) );
  INVX0 U803 ( .INP(G13), .ZN(n776) );
  XNOR2X1 U804 ( .IN1(n781), .IN2(keyinput154), .Q(n779) );
  NAND2X0 U805 ( .IN1(n622), .IN2(n664), .QN(n781) );
  XOR2X1 U806 ( .IN1(n782), .IN2(keyinput143), .Q(n622) );
  NAND2X0 U807 ( .IN1(n704), .IN2(n783), .QN(n782) );
  NOR2X0 U808 ( .IN1(n666), .IN2(n611), .QN(n704) );
  XOR3X1 U809 ( .IN1(keyinput245), .IN2(keyinput227), .IN3(n784), .Q(G1335) );
  NOR2X0 U810 ( .IN1(n785), .IN2(n786), .QN(n784) );
  XOR2X1 U811 ( .IN1(keyinput197), .IN2(n787), .Q(n786) );
  AND2X1 U812 ( .IN1(n788), .IN2(G12), .Q(n787) );
  XOR2X1 U813 ( .IN1(n789), .IN2(keyinput198), .Q(n785) );
  NAND2X0 U814 ( .IN1(n788), .IN2(n790), .QN(n789) );
  XNOR2X1 U815 ( .IN1(n791), .IN2(keyinput172), .Q(n788) );
  NAND2X0 U816 ( .IN1(G12), .IN2(n790), .QN(n791) );
  XNOR2X1 U817 ( .IN1(n792), .IN2(keyinput153), .Q(n790) );
  NAND2X0 U818 ( .IN1(n634), .IN2(n623), .QN(n792) );
  XOR3X1 U819 ( .IN1(keyinput243), .IN2(keyinput225), .IN3(n793), .Q(G1333) );
  NOR2X0 U820 ( .IN1(n794), .IN2(n795), .QN(n793) );
  XOR2X1 U821 ( .IN1(keyinput193), .IN2(n796), .Q(n795) );
  NOR2X0 U822 ( .IN1(n797), .IN2(n798), .QN(n796) );
  XOR2X1 U823 ( .IN1(keyinput194), .IN2(n799), .Q(n794) );
  NOR2X0 U824 ( .IN1(n800), .IN2(n798), .QN(n799) );
  XNOR2X1 U825 ( .IN1(n801), .IN2(keyinput170), .Q(n798) );
  OR2X1 U826 ( .IN1(n797), .IN2(n800), .Q(n801) );
  XOR2X1 U827 ( .IN1(n802), .IN2(keyinput151), .Q(n800) );
  NAND2X0 U828 ( .IN1(n634), .IN2(n680), .QN(n802) );
  XOR3X1 U829 ( .IN1(keyinput242), .IN2(keyinput224), .IN3(n803), .Q(G1332) );
  NOR2X0 U830 ( .IN1(n804), .IN2(n805), .QN(n803) );
  XOR2X1 U831 ( .IN1(keyinput191), .IN2(n806), .Q(n805) );
  NOR2X0 U832 ( .IN1(n807), .IN2(n808), .QN(n806) );
  XOR2X1 U833 ( .IN1(keyinput192), .IN2(n809), .Q(n804) );
  NOR2X0 U834 ( .IN1(n807), .IN2(n810), .QN(n809) );
  XOR2X1 U835 ( .IN1(n811), .IN2(keyinput169), .Q(n807) );
  OR2X1 U836 ( .IN1(n810), .IN2(n808), .Q(n811) );
  XNOR2X1 U837 ( .IN1(n812), .IN2(keyinput150), .Q(n810) );
  NAND2X0 U838 ( .IN1(n634), .IN2(n664), .QN(n812) );
  XOR2X1 U839 ( .IN1(n813), .IN2(keyinput142), .Q(n634) );
  NAND3X0 U840 ( .IN1(n611), .IN2(n666), .IN3(n783), .QN(n813) );
  AND3X1 U841 ( .IN1(n814), .IN2(n690), .IN3(n675), .Q(n783) );
  INVX0 U842 ( .INP(n677), .ZN(n690) );
  XOR3X1 U843 ( .IN1(keyinput239), .IN2(keyinput221), .IN3(n815), .Q(G1325) );
  NOR2X0 U844 ( .IN1(n816), .IN2(n817), .QN(n815) );
  XOR2X1 U845 ( .IN1(keyinput185), .IN2(n818), .Q(n817) );
  NOR2X0 U846 ( .IN1(n819), .IN2(n820), .QN(n818) );
  XOR2X1 U847 ( .IN1(keyinput186), .IN2(n821), .Q(n816) );
  NOR2X0 U848 ( .IN1(n822), .IN2(n820), .QN(n821) );
  XNOR2X1 U849 ( .IN1(n823), .IN2(keyinput166), .Q(n820) );
  OR2X1 U850 ( .IN1(n822), .IN2(n819), .Q(n823) );
  XNOR2X1 U851 ( .IN1(n824), .IN2(keyinput147), .Q(n822) );
  NAND2X0 U852 ( .IN1(n645), .IN2(n680), .QN(n824) );
  XOR2X1 U853 ( .IN1(n825), .IN2(keyinput141), .Q(n645) );
  NAND3X0 U854 ( .IN1(n611), .IN2(n666), .IN3(n703), .QN(n825) );
  AND3X1 U855 ( .IN1(n814), .IN2(n687), .IN3(n677), .Q(n703) );
  MUX21X1 U856 ( .IN1(n826), .IN2(n827), .S(n828), .Q(n677) );
  XOR3X1 U857 ( .IN1(G21), .IN2(G17), .IN3(n829), .Q(n828) );
  XOR2X1 U858 ( .IN1(G29), .IN2(G25), .Q(n829) );
  NAND2X0 U859 ( .IN1(n830), .IN2(n831), .QN(n827) );
  AND2X1 U860 ( .IN1(n831), .IN2(n830), .Q(n826) );
  NAND3X0 U861 ( .IN1(G41), .IN2(n832), .IN3(G37), .QN(n830) );
  AO21X1 U862 ( .IN1(G37), .IN2(G41), .IN3(n832), .Q(n831) );
  XOR2X1 U863 ( .IN1(n833), .IN2(n834), .Q(n832) );
  INVX0 U864 ( .INP(n675), .ZN(n687) );
  MUX21X1 U865 ( .IN1(n835), .IN2(n836), .S(n837), .Q(n675) );
  XOR3X1 U866 ( .IN1(G22), .IN2(G18), .IN3(n838), .Q(n837) );
  XOR2X1 U867 ( .IN1(G30), .IN2(G26), .Q(n838) );
  NAND2X0 U868 ( .IN1(n839), .IN2(n840), .QN(n836) );
  AND2X1 U869 ( .IN1(n840), .IN2(n839), .Q(n835) );
  NAND3X0 U870 ( .IN1(G41), .IN2(n841), .IN3(G38), .QN(n839) );
  AO21X1 U871 ( .IN1(G38), .IN2(G41), .IN3(n841), .Q(n840) );
  XOR2X1 U872 ( .IN1(n842), .IN2(n843), .Q(n841) );
  XNOR2X1 U873 ( .IN1(n844), .IN2(keyinput140), .Q(n814) );
  NAND3X0 U874 ( .IN1(n845), .IN2(n846), .IN3(n847), .QN(n844) );
  OA222X1 U875 ( .IN1(n848), .IN2(n849), .IN3(n850), .IN4(n851), .IN5(n852), 
        .IN6(n853), .Q(n847) );
  INVX0 U876 ( .INP(keyinput137), .ZN(n853) );
  NOR2X0 U877 ( .IN1(n849), .IN2(n635), .QN(n852) );
  INVX0 U878 ( .INP(keyinput136), .ZN(n851) );
  NOR2X0 U879 ( .IN1(n680), .IN2(n849), .QN(n850) );
  INVX0 U880 ( .INP(n691), .ZN(n849) );
  NOR2X0 U881 ( .IN1(n623), .IN2(n664), .QN(n691) );
  OA22X1 U882 ( .IN1(keyinput137), .IN2(n635), .IN3(keyinput136), .IN4(n680), 
        .Q(n848) );
  XOR2X1 U883 ( .IN1(keyinput138), .IN2(n854), .Q(n846) );
  NOR2X0 U884 ( .IN1(n623), .IN2(n855), .QN(n854) );
  XOR2X1 U885 ( .IN1(n856), .IN2(keyinput132), .Q(n623) );
  NAND2X0 U886 ( .IN1(n857), .IN2(n858), .QN(n856) );
  XOR2X1 U887 ( .IN1(n859), .IN2(keyinput128), .Q(n858) );
  NAND2X0 U888 ( .IN1(n860), .IN2(n861), .QN(n859) );
  XOR2X1 U889 ( .IN1(n862), .IN2(keyinput127), .Q(n857) );
  NAND2X0 U890 ( .IN1(n860), .IN2(n863), .QN(n862) );
  XNOR2X1 U891 ( .IN1(n864), .IN2(keyinput120), .Q(n860) );
  NAND2X0 U892 ( .IN1(n863), .IN2(n861), .QN(n864) );
  XNOR2X1 U893 ( .IN1(n865), .IN2(keyinput116), .Q(n861) );
  NAND2X0 U894 ( .IN1(n866), .IN2(n867), .QN(n865) );
  XOR2X1 U895 ( .IN1(keyinput112), .IN2(n868), .Q(n867) );
  NOR2X0 U896 ( .IN1(n869), .IN2(n870), .QN(n868) );
  XOR2X1 U897 ( .IN1(keyinput100), .IN2(n871), .Q(n870) );
  XOR2X1 U898 ( .IN1(n872), .IN2(keyinput111), .Q(n866) );
  NAND2X0 U899 ( .IN1(n873), .IN2(n874), .QN(n872) );
  INVX0 U900 ( .INP(n869), .ZN(n873) );
  XOR2X1 U901 ( .IN1(n875), .IN2(keyinput104), .Q(n869) );
  NAND2X0 U902 ( .IN1(n876), .IN2(n874), .QN(n875) );
  XNOR2X1 U903 ( .IN1(n877), .IN2(keyinput3), .Q(n874) );
  NAND2X0 U904 ( .IN1(G36), .IN2(G41), .QN(n877) );
  XNOR2X1 U905 ( .IN1(keyinput100), .IN2(n871), .Q(n876) );
  AND2X1 U906 ( .IN1(n878), .IN2(n879), .Q(n871) );
  XOR2X1 U907 ( .IN1(keyinput96), .IN2(n880), .Q(n879) );
  AND2X1 U908 ( .IN1(n881), .IN2(n882), .Q(n880) );
  XOR2X1 U909 ( .IN1(n883), .IN2(keyinput95), .Q(n878) );
  NAND2X0 U910 ( .IN1(n884), .IN2(n882), .QN(n883) );
  XNOR2X1 U911 ( .IN1(n885), .IN2(keyinput88), .Q(n882) );
  NAND2X0 U912 ( .IN1(n884), .IN2(n881), .QN(n885) );
  XNOR2X1 U913 ( .IN1(n886), .IN2(keyinput84), .Q(n863) );
  NAND2X0 U914 ( .IN1(n887), .IN2(n888), .QN(n886) );
  XOR2X1 U915 ( .IN1(n889), .IN2(keyinput76), .Q(n888) );
  NAND2X0 U916 ( .IN1(n890), .IN2(n891), .QN(n889) );
  XOR2X1 U917 ( .IN1(n892), .IN2(keyinput75), .Q(n887) );
  NAND2X0 U918 ( .IN1(n890), .IN2(n893), .QN(n892) );
  XOR2X1 U919 ( .IN1(n894), .IN2(keyinput63), .Q(n890) );
  NAND2X0 U920 ( .IN1(n893), .IN2(n891), .QN(n894) );
  XOR2X1 U921 ( .IN1(n895), .IN2(keyinput55), .Q(n891) );
  NAND2X0 U922 ( .IN1(n896), .IN2(n897), .QN(n895) );
  XOR2X1 U923 ( .IN1(keyinput41), .IN2(n898), .Q(n897) );
  NOR2X0 U924 ( .IN1(n899), .IN2(n900), .QN(n898) );
  XOR2X1 U925 ( .IN1(keyinput42), .IN2(n901), .Q(n896) );
  NOR2X0 U926 ( .IN1(n617), .IN2(n900), .QN(n901) );
  XNOR2X1 U927 ( .IN1(n902), .IN2(keyinput15), .Q(n900) );
  NAND2X0 U928 ( .IN1(G12), .IN2(G16), .QN(n902) );
  INVX0 U929 ( .INP(G16), .ZN(n617) );
  XOR2X1 U930 ( .IN1(n903), .IN2(keyinput54), .Q(n893) );
  NAND2X0 U931 ( .IN1(n904), .IN2(n905), .QN(n903) );
  XOR2X1 U932 ( .IN1(n906), .IN2(keyinput39), .Q(n905) );
  NAND2X0 U933 ( .IN1(G4), .IN2(n907), .QN(n906) );
  XOR2X1 U934 ( .IN1(n908), .IN2(keyinput40), .Q(n904) );
  NAND2X0 U935 ( .IN1(G8), .IN2(n907), .QN(n908) );
  XNOR2X1 U936 ( .IN1(n909), .IN2(keyinput14), .Q(n907) );
  NAND2X0 U937 ( .IN1(G4), .IN2(G8), .QN(n909) );
  MUX21X1 U938 ( .IN1(n910), .IN2(n911), .S(keyinput135), .Q(n845) );
  OR2X1 U939 ( .IN1(n855), .IN2(n664), .Q(n911) );
  NOR2X0 U940 ( .IN1(n664), .IN2(n855), .QN(n910) );
  INVX0 U941 ( .INP(n727), .ZN(n855) );
  NOR2X0 U942 ( .IN1(n635), .IN2(n680), .QN(n727) );
  XOR2X1 U943 ( .IN1(n912), .IN2(keyinput130), .Q(n680) );
  NAND2X0 U944 ( .IN1(n913), .IN2(n914), .QN(n912) );
  XOR2X1 U945 ( .IN1(keyinput123), .IN2(n915), .Q(n914) );
  NOR2X0 U946 ( .IN1(n916), .IN2(n917), .QN(n915) );
  INVX0 U947 ( .INP(n918), .ZN(n917) );
  XOR2X1 U948 ( .IN1(n919), .IN2(keyinput82), .Q(n916) );
  XOR2X1 U949 ( .IN1(n920), .IN2(keyinput124), .Q(n913) );
  NAND2X0 U950 ( .IN1(n918), .IN2(n921), .QN(n920) );
  XOR2X1 U951 ( .IN1(n922), .IN2(keyinput118), .Q(n918) );
  NAND2X0 U952 ( .IN1(n921), .IN2(n923), .QN(n922) );
  XNOR2X1 U953 ( .IN1(keyinput82), .IN2(n919), .Q(n923) );
  AO21X1 U954 ( .IN1(n924), .IN2(n925), .IN3(n926), .Q(n919) );
  XOR2X1 U955 ( .IN1(n927), .IN2(keyinput72), .Q(n926) );
  NAND3X0 U956 ( .IN1(n928), .IN2(n929), .IN3(n930), .QN(n927) );
  INVX0 U957 ( .INP(keyinput61), .ZN(n929) );
  XOR2X1 U958 ( .IN1(n928), .IN2(keyinput61), .Q(n924) );
  NAND2X0 U959 ( .IN1(n930), .IN2(n925), .QN(n928) );
  XOR2X1 U960 ( .IN1(G10), .IN2(G14), .Q(n925) );
  XOR2X1 U961 ( .IN1(keyinput51), .IN2(n931), .Q(n930) );
  OA21X1 U962 ( .IN1(G6), .IN2(n819), .IN3(n932), .Q(n931) );
  XOR2X1 U963 ( .IN1(keyinput34), .IN2(n933), .Q(n932) );
  AND2X1 U964 ( .IN1(n819), .IN2(G6), .Q(n933) );
  INVX0 U965 ( .INP(G2), .ZN(n819) );
  XOR2X1 U966 ( .IN1(n934), .IN2(keyinput114), .Q(n921) );
  NAND2X0 U967 ( .IN1(n935), .IN2(n936), .QN(n934) );
  XOR2X1 U968 ( .IN1(n937), .IN2(keyinput108), .Q(n936) );
  NAND2X0 U969 ( .IN1(n938), .IN2(n939), .QN(n937) );
  XOR2X1 U970 ( .IN1(n940), .IN2(keyinput107), .Q(n935) );
  NAND2X0 U971 ( .IN1(n941), .IN2(n939), .QN(n940) );
  XNOR2X1 U972 ( .IN1(n942), .IN2(keyinput102), .Q(n939) );
  NAND2X0 U973 ( .IN1(n938), .IN2(n941), .QN(n942) );
  XOR2X1 U974 ( .IN1(n943), .IN2(keyinput98), .Q(n938) );
  NAND2X0 U975 ( .IN1(n944), .IN2(n945), .QN(n943) );
  XOR2X1 U976 ( .IN1(keyinput91), .IN2(n946), .Q(n945) );
  NOR2X0 U977 ( .IN1(n947), .IN2(n948), .QN(n946) );
  XOR2X1 U978 ( .IN1(keyinput92), .IN2(n949), .Q(n944) );
  NOR2X0 U979 ( .IN1(n950), .IN2(n948), .QN(n949) );
  XNOR2X1 U980 ( .IN1(n951), .IN2(keyinput86), .Q(n948) );
  NAND2X0 U981 ( .IN1(n952), .IN2(n881), .QN(n951) );
  INVX0 U982 ( .INP(n950), .ZN(n881) );
  XOR2X1 U983 ( .IN1(n953), .IN2(keyinput81), .Q(n950) );
  NAND2X0 U984 ( .IN1(n954), .IN2(n955), .QN(n953) );
  XOR2X1 U985 ( .IN1(keyinput70), .IN2(n956), .Q(n955) );
  NOR2X0 U986 ( .IN1(n957), .IN2(n958), .QN(n956) );
  XNOR2X1 U987 ( .IN1(keyinput49), .IN2(n959), .Q(n958) );
  XOR2X1 U988 ( .IN1(keyinput71), .IN2(n960), .Q(n954) );
  NOR2X0 U989 ( .IN1(n957), .IN2(n961), .QN(n960) );
  XNOR2X1 U990 ( .IN1(keyinput50), .IN2(n962), .Q(n961) );
  XNOR2X1 U991 ( .IN1(n963), .IN2(keyinput60), .Q(n957) );
  NAND2X0 U992 ( .IN1(n964), .IN2(n965), .QN(n963) );
  XOR2X1 U993 ( .IN1(n959), .IN2(keyinput49), .Q(n965) );
  NAND2X0 U994 ( .IN1(n966), .IN2(n967), .QN(n959) );
  XOR2X1 U995 ( .IN1(keyinput30), .IN2(n968), .Q(n967) );
  AND2X1 U996 ( .IN1(n969), .IN2(G29), .Q(n968) );
  XOR2X1 U997 ( .IN1(n970), .IN2(keyinput31), .Q(n966) );
  NAND2X0 U998 ( .IN1(G30), .IN2(n969), .QN(n970) );
  XNOR2X1 U999 ( .IN1(n971), .IN2(keyinput10), .Q(n969) );
  NAND2X0 U1000 ( .IN1(G29), .IN2(G30), .QN(n971) );
  XOR2X1 U1001 ( .IN1(n962), .IN2(keyinput50), .Q(n964) );
  NAND2X0 U1002 ( .IN1(n972), .IN2(n973), .QN(n962) );
  XOR2X1 U1003 ( .IN1(keyinput32), .IN2(n974), .Q(n973) );
  NOR2X0 U1004 ( .IN1(n975), .IN2(n671), .QN(n974) );
  INVX0 U1005 ( .INP(G31), .ZN(n671) );
  XOR2X1 U1006 ( .IN1(keyinput33), .IN2(n976), .Q(n972) );
  NOR2X0 U1007 ( .IN1(n975), .IN2(n977), .QN(n976) );
  INVX0 U1008 ( .INP(G32), .ZN(n977) );
  XOR2X1 U1009 ( .IN1(n978), .IN2(keyinput11), .Q(n975) );
  NAND2X0 U1010 ( .IN1(G31), .IN2(G32), .QN(n978) );
  XOR2X1 U1011 ( .IN1(n979), .IN2(keyinput1), .Q(n941) );
  NAND2X0 U1012 ( .IN1(G34), .IN2(G41), .QN(n979) );
  INVX0 U1013 ( .INP(n678), .ZN(n635) );
  XOR2X1 U1014 ( .IN1(n980), .IN2(keyinput131), .Q(n678) );
  NAND2X0 U1015 ( .IN1(n981), .IN2(n982), .QN(n980) );
  XOR2X1 U1016 ( .IN1(keyinput125), .IN2(n983), .Q(n982) );
  NOR2X0 U1017 ( .IN1(n984), .IN2(n985), .QN(n983) );
  XNOR2X1 U1018 ( .IN1(keyinput83), .IN2(n986), .Q(n985) );
  XOR2X1 U1019 ( .IN1(n987), .IN2(keyinput126), .Q(n981) );
  NAND2X0 U1020 ( .IN1(n988), .IN2(n989), .QN(n987) );
  INVX0 U1021 ( .INP(n984), .ZN(n988) );
  XOR2X1 U1022 ( .IN1(n990), .IN2(keyinput119), .Q(n984) );
  NAND2X0 U1023 ( .IN1(n991), .IN2(n989), .QN(n990) );
  XNOR2X1 U1024 ( .IN1(n992), .IN2(keyinput115), .Q(n989) );
  NAND2X0 U1025 ( .IN1(n993), .IN2(n994), .QN(n992) );
  XOR2X1 U1026 ( .IN1(keyinput109), .IN2(n995), .Q(n994) );
  NOR2X0 U1027 ( .IN1(n996), .IN2(n997), .QN(n995) );
  XNOR2X1 U1028 ( .IN1(keyinput103), .IN2(n998), .Q(n997) );
  XOR2X1 U1029 ( .IN1(n999), .IN2(keyinput110), .Q(n993) );
  NAND2X0 U1030 ( .IN1(n1000), .IN2(n1001), .QN(n999) );
  XOR2X1 U1031 ( .IN1(keyinput103), .IN2(n998), .Q(n1000) );
  NOR2X0 U1032 ( .IN1(n1002), .IN2(n996), .QN(n998) );
  XOR2X1 U1033 ( .IN1(n1003), .IN2(keyinput2), .Q(n996) );
  NAND2X0 U1034 ( .IN1(G35), .IN2(G41), .QN(n1003) );
  INVX0 U1035 ( .INP(n1001), .ZN(n1002) );
  XNOR2X1 U1036 ( .IN1(n1004), .IN2(keyinput99), .Q(n1001) );
  NAND2X0 U1037 ( .IN1(n1005), .IN2(n1006), .QN(n1004) );
  XOR2X1 U1038 ( .IN1(keyinput93), .IN2(n1007), .Q(n1006) );
  NOR2X0 U1039 ( .IN1(n1008), .IN2(n1009), .QN(n1007) );
  XOR2X1 U1040 ( .IN1(n1010), .IN2(keyinput94), .Q(n1005) );
  OR2X1 U1041 ( .IN1(n1009), .IN2(n947), .Q(n1010) );
  INVX0 U1042 ( .INP(n952), .ZN(n947) );
  XNOR2X1 U1043 ( .IN1(n1011), .IN2(keyinput87), .Q(n1009) );
  NAND2X0 U1044 ( .IN1(n952), .IN2(n1012), .QN(n1011) );
  XOR2X1 U1045 ( .IN1(n1013), .IN2(keyinput80), .Q(n952) );
  NAND2X0 U1046 ( .IN1(n1014), .IN2(n1015), .QN(n1013) );
  XOR2X1 U1047 ( .IN1(keyinput68), .IN2(n1016), .Q(n1015) );
  NOR2X0 U1048 ( .IN1(n1017), .IN2(n1018), .QN(n1016) );
  XOR2X1 U1049 ( .IN1(keyinput47), .IN2(n1019), .Q(n1018) );
  XOR2X1 U1050 ( .IN1(keyinput69), .IN2(n1020), .Q(n1014) );
  NOR2X0 U1051 ( .IN1(n1021), .IN2(n1017), .QN(n1020) );
  XNOR2X1 U1052 ( .IN1(n1022), .IN2(keyinput59), .Q(n1017) );
  NAND2X0 U1053 ( .IN1(n1023), .IN2(n1024), .QN(n1022) );
  XNOR2X1 U1054 ( .IN1(keyinput48), .IN2(n1025), .Q(n1024) );
  XNOR2X1 U1055 ( .IN1(keyinput47), .IN2(n1019), .Q(n1023) );
  AND2X1 U1056 ( .IN1(n1026), .IN2(n1027), .Q(n1019) );
  XOR2X1 U1057 ( .IN1(keyinput26), .IN2(n1028), .Q(n1027) );
  NOR2X0 U1058 ( .IN1(n688), .IN2(n1029), .QN(n1028) );
  INVX0 U1059 ( .INP(G25), .ZN(n688) );
  XOR2X1 U1060 ( .IN1(keyinput27), .IN2(n1030), .Q(n1026) );
  NOR2X0 U1061 ( .IN1(n685), .IN2(n1029), .QN(n1030) );
  XNOR2X1 U1062 ( .IN1(n1031), .IN2(keyinput8), .Q(n1029) );
  NAND2X0 U1063 ( .IN1(G25), .IN2(G26), .QN(n1031) );
  INVX0 U1064 ( .INP(G26), .ZN(n685) );
  XOR2X1 U1065 ( .IN1(n1025), .IN2(keyinput48), .Q(n1021) );
  NAND2X0 U1066 ( .IN1(n1032), .IN2(n1033), .QN(n1025) );
  XOR2X1 U1067 ( .IN1(n1034), .IN2(keyinput28), .Q(n1033) );
  NAND2X0 U1068 ( .IN1(n1035), .IN2(G27), .QN(n1034) );
  XOR2X1 U1069 ( .IN1(n1036), .IN2(keyinput29), .Q(n1032) );
  NAND2X0 U1070 ( .IN1(n1035), .IN2(G28), .QN(n1036) );
  XOR2X1 U1071 ( .IN1(n1037), .IN2(keyinput9), .Q(n1035) );
  NAND2X0 U1072 ( .IN1(G27), .IN2(G28), .QN(n1037) );
  XOR2X1 U1073 ( .IN1(n986), .IN2(keyinput83), .Q(n991) );
  NAND2X0 U1074 ( .IN1(n1038), .IN2(n1039), .QN(n986) );
  XOR2X1 U1075 ( .IN1(keyinput74), .IN2(n1040), .Q(n1039) );
  NOR2X0 U1076 ( .IN1(n1041), .IN2(n1042), .QN(n1040) );
  XOR2X1 U1077 ( .IN1(n1043), .IN2(keyinput53), .Q(n1042) );
  XOR2X1 U1078 ( .IN1(n1044), .IN2(keyinput73), .Q(n1038) );
  NAND2X0 U1079 ( .IN1(n1045), .IN2(n1046), .QN(n1044) );
  INVX0 U1080 ( .INP(n1041), .ZN(n1046) );
  XOR2X1 U1081 ( .IN1(n1047), .IN2(keyinput62), .Q(n1041) );
  NAND2X0 U1082 ( .IN1(n1045), .IN2(n1048), .QN(n1047) );
  XNOR2X1 U1083 ( .IN1(keyinput53), .IN2(n1043), .Q(n1048) );
  NAND2X0 U1084 ( .IN1(n1049), .IN2(n1050), .QN(n1043) );
  XOR2X1 U1085 ( .IN1(n1051), .IN2(keyinput37), .Q(n1050) );
  NAND2X0 U1086 ( .IN1(n1052), .IN2(G11), .QN(n1051) );
  XOR2X1 U1087 ( .IN1(n1053), .IN2(keyinput38), .Q(n1049) );
  NAND2X0 U1088 ( .IN1(n1052), .IN2(G15), .QN(n1053) );
  XOR2X1 U1089 ( .IN1(n1054), .IN2(keyinput13), .Q(n1052) );
  NAND2X0 U1090 ( .IN1(G11), .IN2(G15), .QN(n1054) );
  XOR2X1 U1091 ( .IN1(n1055), .IN2(keyinput52), .Q(n1045) );
  NAND2X0 U1092 ( .IN1(n1056), .IN2(n1057), .QN(n1055) );
  XOR2X1 U1093 ( .IN1(n1058), .IN2(keyinput35), .Q(n1057) );
  NAND2X0 U1094 ( .IN1(G3), .IN2(n1059), .QN(n1058) );
  XOR2X1 U1095 ( .IN1(n1060), .IN2(keyinput36), .Q(n1056) );
  NAND2X0 U1096 ( .IN1(G7), .IN2(n1059), .QN(n1060) );
  XNOR2X1 U1097 ( .IN1(n1061), .IN2(keyinput12), .Q(n1059) );
  NAND2X0 U1098 ( .IN1(G3), .IN2(G7), .QN(n1061) );
  XOR2X1 U1099 ( .IN1(n1062), .IN2(keyinput129), .Q(n664) );
  NAND2X0 U1100 ( .IN1(n1063), .IN2(n1064), .QN(n1062) );
  XOR2X1 U1101 ( .IN1(keyinput121), .IN2(n1065), .Q(n1064) );
  NOR2X0 U1102 ( .IN1(n1066), .IN2(n1067), .QN(n1065) );
  XOR2X1 U1103 ( .IN1(keyinput122), .IN2(n1068), .Q(n1063) );
  NOR2X0 U1104 ( .IN1(n1069), .IN2(n1067), .QN(n1068) );
  XNOR2X1 U1105 ( .IN1(n1070), .IN2(keyinput117), .Q(n1067) );
  NAND2X0 U1106 ( .IN1(n1071), .IN2(n1072), .QN(n1070) );
  INVX0 U1107 ( .INP(n1066), .ZN(n1072) );
  XOR3X1 U1108 ( .IN1(G13), .IN2(G1), .IN3(n1073), .Q(n1066) );
  XOR2X1 U1109 ( .IN1(G5), .IN2(n808), .Q(n1073) );
  INVX0 U1110 ( .INP(G9), .ZN(n808) );
  XNOR2X1 U1111 ( .IN1(keyinput113), .IN2(n1074), .Q(n1071) );
  XOR2X1 U1112 ( .IN1(n1074), .IN2(keyinput113), .Q(n1069) );
  NAND2X0 U1113 ( .IN1(n1075), .IN2(n1076), .QN(n1074) );
  XOR2X1 U1114 ( .IN1(n1077), .IN2(keyinput106), .Q(n1076) );
  NAND2X0 U1115 ( .IN1(n1078), .IN2(n1079), .QN(n1077) );
  XOR2X1 U1116 ( .IN1(n1080), .IN2(keyinput105), .Q(n1075) );
  NAND2X0 U1117 ( .IN1(n1078), .IN2(n1081), .QN(n1080) );
  XNOR2X1 U1118 ( .IN1(n1082), .IN2(keyinput101), .Q(n1078) );
  NAND2X0 U1119 ( .IN1(n1081), .IN2(n1079), .QN(n1082) );
  XNOR2X1 U1120 ( .IN1(n1083), .IN2(keyinput97), .Q(n1079) );
  NAND2X0 U1121 ( .IN1(n1084), .IN2(n1085), .QN(n1083) );
  XOR2X1 U1122 ( .IN1(keyinput89), .IN2(n1086), .Q(n1085) );
  AND2X1 U1123 ( .IN1(n1012), .IN2(n1087), .Q(n1086) );
  XOR2X1 U1124 ( .IN1(n1088), .IN2(keyinput90), .Q(n1084) );
  NAND2X0 U1125 ( .IN1(n884), .IN2(n1087), .QN(n1088) );
  XNOR2X1 U1126 ( .IN1(n1089), .IN2(keyinput85), .Q(n1087) );
  NAND2X0 U1127 ( .IN1(n884), .IN2(n1012), .QN(n1089) );
  INVX0 U1128 ( .INP(n1008), .ZN(n1012) );
  XOR2X1 U1129 ( .IN1(n1090), .IN2(keyinput78), .Q(n1008) );
  NAND2X0 U1130 ( .IN1(n1091), .IN2(n1092), .QN(n1090) );
  XOR2X1 U1131 ( .IN1(keyinput64), .IN2(n1093), .Q(n1092) );
  NOR2X0 U1132 ( .IN1(n1094), .IN2(n1095), .QN(n1093) );
  XOR2X1 U1133 ( .IN1(n1096), .IN2(keyinput43), .Q(n1095) );
  XOR2X1 U1134 ( .IN1(keyinput65), .IN2(n1097), .Q(n1091) );
  NOR2X0 U1135 ( .IN1(n1094), .IN2(n1098), .QN(n1097) );
  XOR2X1 U1136 ( .IN1(keyinput44), .IN2(n1099), .Q(n1098) );
  XOR2X1 U1137 ( .IN1(n1100), .IN2(keyinput57), .Q(n1094) );
  NAND2X0 U1138 ( .IN1(n1101), .IN2(n1102), .QN(n1100) );
  XNOR2X1 U1139 ( .IN1(keyinput43), .IN2(n1096), .Q(n1102) );
  NAND2X0 U1140 ( .IN1(n1103), .IN2(n1104), .QN(n1096) );
  XOR2X1 U1141 ( .IN1(keyinput18), .IN2(n1105), .Q(n1104) );
  AND2X1 U1142 ( .IN1(n1106), .IN2(G17), .Q(n1105) );
  XOR2X1 U1143 ( .IN1(n1107), .IN2(keyinput19), .Q(n1103) );
  NAND2X0 U1144 ( .IN1(G18), .IN2(n1106), .QN(n1107) );
  XNOR2X1 U1145 ( .IN1(n1108), .IN2(keyinput4), .Q(n1106) );
  NAND2X0 U1146 ( .IN1(G17), .IN2(G18), .QN(n1108) );
  XNOR2X1 U1147 ( .IN1(keyinput44), .IN2(n1099), .Q(n1101) );
  AND2X1 U1148 ( .IN1(n1109), .IN2(n1110), .Q(n1099) );
  XOR2X1 U1149 ( .IN1(n1111), .IN2(keyinput20), .Q(n1110) );
  NAND2X0 U1150 ( .IN1(G19), .IN2(n1112), .QN(n1111) );
  XOR2X1 U1151 ( .IN1(n1113), .IN2(keyinput21), .Q(n1109) );
  NAND2X0 U1152 ( .IN1(G20), .IN2(n1112), .QN(n1113) );
  XNOR2X1 U1153 ( .IN1(n1114), .IN2(keyinput5), .Q(n1112) );
  NAND2X0 U1154 ( .IN1(G19), .IN2(G20), .QN(n1114) );
  XOR2X1 U1155 ( .IN1(n1115), .IN2(keyinput79), .Q(n884) );
  NAND2X0 U1156 ( .IN1(n1116), .IN2(n1117), .QN(n1115) );
  XOR2X1 U1157 ( .IN1(keyinput67), .IN2(n1118), .Q(n1117) );
  NOR2X0 U1158 ( .IN1(n1119), .IN2(n1120), .QN(n1118) );
  XOR2X1 U1159 ( .IN1(n1121), .IN2(keyinput46), .Q(n1120) );
  XOR2X1 U1160 ( .IN1(n1122), .IN2(keyinput66), .Q(n1116) );
  NAND2X0 U1161 ( .IN1(n1123), .IN2(n1124), .QN(n1122) );
  INVX0 U1162 ( .INP(n1119), .ZN(n1124) );
  XOR2X1 U1163 ( .IN1(n1125), .IN2(keyinput58), .Q(n1119) );
  NAND2X0 U1164 ( .IN1(n1123), .IN2(n1126), .QN(n1125) );
  XNOR2X1 U1165 ( .IN1(keyinput46), .IN2(n1121), .Q(n1126) );
  NAND2X0 U1166 ( .IN1(n1127), .IN2(n1128), .QN(n1121) );
  XOR2X1 U1167 ( .IN1(keyinput24), .IN2(n1129), .Q(n1128) );
  NOR2X0 U1168 ( .IN1(n693), .IN2(n1130), .QN(n1129) );
  INVX0 U1169 ( .INP(G23), .ZN(n693) );
  XOR2X1 U1170 ( .IN1(n1131), .IN2(keyinput25), .Q(n1127) );
  OR2X1 U1171 ( .IN1(n1130), .IN2(n710), .Q(n1131) );
  INVX0 U1172 ( .INP(G24), .ZN(n710) );
  XNOR2X1 U1173 ( .IN1(n1132), .IN2(keyinput7), .Q(n1130) );
  NAND2X0 U1174 ( .IN1(G23), .IN2(G24), .QN(n1132) );
  XOR2X1 U1175 ( .IN1(n1133), .IN2(keyinput45), .Q(n1123) );
  NAND2X0 U1176 ( .IN1(n1134), .IN2(n1135), .QN(n1133) );
  XOR2X1 U1177 ( .IN1(keyinput22), .IN2(n1136), .Q(n1135) );
  NOR2X0 U1178 ( .IN1(n696), .IN2(n1137), .QN(n1136) );
  INVX0 U1179 ( .INP(G21), .ZN(n696) );
  XOR2X1 U1180 ( .IN1(keyinput23), .IN2(n1138), .Q(n1134) );
  NOR2X0 U1181 ( .IN1(n721), .IN2(n1137), .QN(n1138) );
  XNOR2X1 U1182 ( .IN1(n1139), .IN2(keyinput6), .Q(n1137) );
  NAND2X0 U1183 ( .IN1(G21), .IN2(G22), .QN(n1139) );
  INVX0 U1184 ( .INP(G22), .ZN(n721) );
  XNOR2X1 U1185 ( .IN1(n1140), .IN2(keyinput0), .Q(n1081) );
  NAND2X0 U1186 ( .IN1(G33), .IN2(G41), .QN(n1140) );
  INVX0 U1187 ( .INP(n600), .ZN(n666) );
  MUX21X1 U1188 ( .IN1(n1141), .IN2(n1142), .S(n1143), .Q(n600) );
  XOR3X1 U1189 ( .IN1(G24), .IN2(G20), .IN3(n1144), .Q(n1143) );
  XOR2X1 U1190 ( .IN1(G32), .IN2(G28), .Q(n1144) );
  NAND2X0 U1191 ( .IN1(n1145), .IN2(n1146), .QN(n1142) );
  AND2X1 U1192 ( .IN1(n1146), .IN2(n1145), .Q(n1141) );
  NAND3X0 U1193 ( .IN1(G41), .IN2(G40), .IN3(n1147), .QN(n1145) );
  AO21X1 U1194 ( .IN1(G41), .IN2(G40), .IN3(n1147), .Q(n1146) );
  XNOR2X1 U1195 ( .IN1(n842), .IN2(n833), .Q(n1147) );
  XOR3X1 U1196 ( .IN1(G6), .IN2(n1148), .IN3(G5), .Q(n833) );
  OA21X1 U1197 ( .IN1(G8), .IN2(n1149), .IN3(n1150), .Q(n1148) );
  XOR2X1 U1198 ( .IN1(n1151), .IN2(keyinput17), .Q(n1150) );
  NAND2X0 U1199 ( .IN1(G8), .IN2(n1149), .QN(n1151) );
  INVX0 U1200 ( .INP(G7), .ZN(n1149) );
  XOR2X1 U1201 ( .IN1(keyinput77), .IN2(n1152), .Q(n842) );
  OA21X1 U1202 ( .IN1(n1153), .IN2(n1154), .IN3(n1155), .Q(n1152) );
  XOR2X1 U1203 ( .IN1(n1156), .IN2(keyinput56), .Q(n1155) );
  NAND2X0 U1204 ( .IN1(n1154), .IN2(n1153), .QN(n1156) );
  XOR2X1 U1205 ( .IN1(G16), .IN2(G15), .Q(n1154) );
  XOR2X1 U1206 ( .IN1(G14), .IN2(G13), .Q(n1153) );
  MUX21X1 U1207 ( .IN1(n1157), .IN2(n1158), .S(n1159), .Q(n611) );
  XOR3X1 U1208 ( .IN1(G23), .IN2(G19), .IN3(n1160), .Q(n1159) );
  XOR2X1 U1209 ( .IN1(G31), .IN2(G27), .Q(n1160) );
  NAND2X0 U1210 ( .IN1(n1161), .IN2(n1162), .QN(n1158) );
  AND2X1 U1211 ( .IN1(n1162), .IN2(n1161), .Q(n1157) );
  NAND3X0 U1212 ( .IN1(G39), .IN2(G41), .IN3(n1163), .QN(n1161) );
  AO21X1 U1213 ( .IN1(G39), .IN2(G41), .IN3(n1163), .Q(n1162) );
  XNOR2X1 U1214 ( .IN1(n843), .IN2(n834), .Q(n1163) );
  XOR3X1 U1215 ( .IN1(G2), .IN2(n1164), .IN3(G1), .Q(n834) );
  OA21X1 U1216 ( .IN1(G3), .IN2(n1165), .IN3(n1166), .Q(n1164) );
  XOR2X1 U1217 ( .IN1(n1167), .IN2(keyinput16), .Q(n1166) );
  NAND2X0 U1218 ( .IN1(G3), .IN2(n1165), .QN(n1167) );
  INVX0 U1219 ( .INP(G4), .ZN(n1165) );
  XOR3X1 U1220 ( .IN1(G11), .IN2(n797), .IN3(n1168), .Q(n843) );
  XOR2X1 U1221 ( .IN1(n899), .IN2(G9), .Q(n1168) );
  INVX0 U1222 ( .INP(G12), .ZN(n899) );
  INVX0 U1223 ( .INP(G10), .ZN(n797) );
endmodule

