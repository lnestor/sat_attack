
module c5315 ( N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, 
        N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, 
        N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, 
        N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, 
        N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, 
        N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, 
        N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, 
        N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, 
        N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, 
        N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, 
        N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, 
        N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, 
        N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, 
        N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, 
        N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, 
        N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, 
        N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, 
        N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, 
        N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, 
        N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, 
        N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, 
        N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, 
        N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, 
        N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, 
        N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, 
        N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, 
        N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128, keyinput0, 
        keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, 
        keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, 
        keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, 
        keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, 
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, 
        keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, 
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, 
        keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, 
        keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, 
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, 
        keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, 
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, 
        keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, 
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, 
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, 
        keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, 
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, 
        keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, 
        keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, 
        keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, 
        keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, 
        keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, 
        keyinput127 );
  input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37,
         N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79,
         N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106,
         N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136,
         N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164,
         N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197,
         N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234,
         N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273,
         N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315,
         N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358,
         N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422,
         N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545,
         N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583,
         N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610,
         N613, N616, N619, N625, N631, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060,
         N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357,
         N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737,
         N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716,
         N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449,
         N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476,
         N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520,
         N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607,
         N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706,
         N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754,
         N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123,
         N8124, N8127, N8128;
  wire   N1, N137, N141, N293, N299, N549, N592, N1137, N1141, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516;
  assign N3360 = N1;
  assign N3359 = N1;
  assign N3358 = N1;
  assign N3357 = N1;
  assign N2309 = N1;
  assign N2139 = N137;
  assign N2142 = N141;
  assign N709 = N141;
  assign N816 = N293;
  assign N3604 = N299;
  assign N2527 = N299;
  assign N2387 = N549;
  assign N1066 = N592;
  assign N1143 = N1137;
  assign N1142 = N1137;
  assign N2584 = N1141;

  NAND2X0 U897 ( .IN1(n828), .IN2(N137), .QN(N8128) );
  MUX41X1 U898 ( .IN1(n829), .IN3(n830), .IN2(N179), .IN4(N176), .S0(n831), 
        .S1(N580), .Q(n828) );
  NAND2X0 U899 ( .IN1(n832), .IN2(N137), .QN(N8127) );
  MUX21X1 U900 ( .IN1(n833), .IN2(n834), .S(keyinput23), .Q(n832) );
  OA21X1 U901 ( .IN1(N176), .IN2(n835), .IN3(n836), .Q(n834) );
  MUX21X1 U902 ( .IN1(n837), .IN2(n838), .S(n839), .Q(n836) );
  MUX21X1 U903 ( .IN1(n829), .IN2(n830), .S(n840), .Q(n838) );
  OR2X1 U904 ( .IN1(n840), .IN2(N179), .Q(n837) );
  NAND2X0 U905 ( .IN1(N176), .IN2(n841), .QN(n833) );
  AO221X1 U906 ( .IN1(n842), .IN2(n830), .IN3(n843), .IN4(n829), .IN5(n844), 
        .Q(N8124) );
  AO22X1 U907 ( .IN1(N64), .IN2(n845), .IN3(N14), .IN4(n846), .Q(n844) );
  AO221X1 U908 ( .IN1(n847), .IN2(n830), .IN3(n848), .IN4(n829), .IN5(n849), 
        .Q(N8123) );
  AO22X1 U909 ( .IN1(n850), .IN2(N64), .IN3(n851), .IN4(N14), .Q(n849) );
  AO222X1 U910 ( .IN1(n852), .IN2(n853), .IN3(n854), .IN4(n855), .IN5(N97), 
        .IN6(N625), .Q(n829) );
  XNOR2X1 U911 ( .IN1(keyinput105), .IN2(n856), .Q(n854) );
  AO222X1 U912 ( .IN1(n857), .IN2(n855), .IN3(n852), .IN4(n858), .IN5(N94), 
        .IN6(N625), .Q(n830) );
  INVX0 U913 ( .INP(n859), .ZN(n857) );
  AO222X1 U914 ( .IN1(N619), .IN2(n860), .IN3(n855), .IN4(n861), .IN5(N118), 
        .IN6(N625), .Q(N8076) );
  XOR2X1 U915 ( .IN1(keyinput105), .IN2(n856), .Q(n861) );
  AOI22X1 U916 ( .IN1(n862), .IN2(n863), .IN3(n864), .IN4(n865), .QN(n856) );
  OR2X1 U917 ( .IN1(n866), .IN2(n867), .Q(n865) );
  XNOR2X1 U918 ( .IN1(keyinput96), .IN2(n863), .Q(n864) );
  XOR3X1 U919 ( .IN1(n868), .IN2(n869), .IN3(n870), .Q(n863) );
  XNOR2X1 U920 ( .IN1(keyinput63), .IN2(n871), .Q(n870) );
  OA21X1 U921 ( .IN1(N400), .IN2(n872), .IN3(n873), .Q(n871) );
  XOR2X1 U922 ( .IN1(keyinput25), .IN2(n874), .Q(n873) );
  NOR2X0 U923 ( .IN1(n875), .IN2(n876), .QN(n874) );
  MUX21X1 U924 ( .IN1(n877), .IN2(n878), .S(n879), .Q(n876) );
  MUX21X1 U925 ( .IN1(N242), .IN2(N254), .S(n879), .Q(n872) );
  XOR3X1 U926 ( .IN1(n880), .IN2(n881), .IN3(n882), .Q(n869) );
  MUX41X1 U927 ( .IN1(N254), .IN3(n883), .IN2(N242), .IN4(n884), .S0(N389), 
        .S1(N257), .Q(n882) );
  OA21X1 U928 ( .IN1(n878), .IN2(n885), .IN3(n877), .Q(n884) );
  NAND2X0 U929 ( .IN1(N251), .IN2(n885), .QN(n883) );
  INVX0 U930 ( .INP(keyinput12), .ZN(n885) );
  MUX41X1 U931 ( .IN1(N242), .IN3(n877), .IN2(N254), .IN4(n878), .S0(N411), 
        .S1(n886), .Q(n881) );
  MUX41X1 U932 ( .IN1(n887), .IN3(N248), .IN2(n888), .IN4(N251), .S0(N374), 
        .S1(n889), .Q(n880) );
  OA21X1 U933 ( .IN1(N435), .IN2(n890), .IN3(n891), .Q(n868) );
  XOR2X1 U934 ( .IN1(n892), .IN2(keyinput29), .Q(n891) );
  NAND2X0 U935 ( .IN1(n893), .IN2(N435), .QN(n892) );
  MUX21X1 U936 ( .IN1(N248), .IN2(N251), .S(n894), .Q(n893) );
  MUX21X1 U937 ( .IN1(N242), .IN2(N254), .S(n894), .Q(n890) );
  NOR2X0 U938 ( .IN1(n867), .IN2(n866), .QN(n862) );
  XNOR2X1 U939 ( .IN1(n895), .IN2(keyinput91), .Q(n866) );
  NAND2X0 U940 ( .IN1(n896), .IN2(n897), .QN(n895) );
  NOR2X0 U941 ( .IN1(n897), .IN2(n896), .QN(n867) );
  XNOR3X1 U942 ( .IN1(keyinput44), .IN2(n898), .IN3(n899), .Q(n896) );
  MUX41X1 U943 ( .IN1(N254), .IN3(n878), .IN2(N242), .IN4(n877), .S0(N422), 
        .S1(N226), .Q(n899) );
  MUX41X1 U944 ( .IN1(n887), .IN3(N248), .IN2(n888), .IN4(N251), .S0(N468), 
        .S1(n900), .Q(n898) );
  XOR2X1 U945 ( .IN1(n901), .IN2(n902), .Q(n897) );
  MUX21X1 U946 ( .IN1(n903), .IN2(n904), .S(N457), .Q(n901) );
  MUX21X1 U947 ( .IN1(n878), .IN2(n877), .S(N210), .Q(n904) );
  MUX21X1 U948 ( .IN1(n905), .IN2(n906), .S(keyinput21), .Q(n903) );
  MUX21X1 U949 ( .IN1(N254), .IN2(N242), .S(N210), .Q(n906) );
  OR2X1 U950 ( .IN1(n888), .IN2(N210), .Q(n905) );
  NAND2X0 U951 ( .IN1(n853), .IN2(n907), .QN(n860) );
  XOR2X1 U952 ( .IN1(n908), .IN2(n909), .Q(n853) );
  MUX21X1 U953 ( .IN1(n910), .IN2(n911), .S(N566), .Q(n909) );
  XNOR3X1 U954 ( .IN1(n912), .IN2(n913), .IN3(n914), .Q(n911) );
  XOR2X1 U955 ( .IN1(n915), .IN2(n916), .Q(n914) );
  XNOR3X1 U956 ( .IN1(n917), .IN2(n918), .IN3(n919), .Q(n916) );
  XOR2X1 U957 ( .IN1(keyinput125), .IN2(n920), .Q(n919) );
  OA21X1 U958 ( .IN1(n921), .IN2(n922), .IN3(n923), .Q(n920) );
  XOR3X1 U959 ( .IN1(n924), .IN2(n925), .IN3(n926), .Q(n915) );
  XNOR2X1 U960 ( .IN1(n927), .IN2(n928), .Q(n926) );
  OA21X1 U961 ( .IN1(n927), .IN2(n913), .IN3(n929), .Q(n928) );
  NOR2X0 U962 ( .IN1(n930), .IN2(n931), .QN(n927) );
  OR2X1 U963 ( .IN1(n932), .IN2(N374), .Q(n925) );
  NAND2X0 U964 ( .IN1(keyinput123), .IN2(n933), .QN(n924) );
  XNOR3X1 U965 ( .IN1(n934), .IN2(n912), .IN3(n933), .Q(n910) );
  OA21X1 U966 ( .IN1(n935), .IN2(n936), .IN3(n937), .Q(n934) );
  MUX21X1 U967 ( .IN1(n938), .IN2(n921), .S(n939), .Q(n937) );
  NAND2X0 U968 ( .IN1(n935), .IN2(n917), .QN(n938) );
  XNOR2X1 U969 ( .IN1(n939), .IN2(n940), .Q(n936) );
  XNOR2X1 U970 ( .IN1(n941), .IN2(n942), .Q(n939) );
  OA21X1 U971 ( .IN1(n923), .IN2(n943), .IN3(n944), .Q(n942) );
  XOR2X1 U972 ( .IN1(keyinput112), .IN2(n945), .Q(n944) );
  NOR2X0 U973 ( .IN1(n946), .IN2(n947), .QN(n945) );
  XNOR2X1 U974 ( .IN1(n948), .IN2(n949), .Q(n947) );
  INVX0 U975 ( .INP(n923), .ZN(n946) );
  XNOR2X1 U976 ( .IN1(n948), .IN2(n930), .Q(n943) );
  AO21X1 U977 ( .IN1(n950), .IN2(n951), .IN3(keyinput94), .Q(n948) );
  OR2X1 U978 ( .IN1(n952), .IN2(n913), .Q(n951) );
  XNOR2X1 U979 ( .IN1(n953), .IN2(n954), .Q(n950) );
  OA21X1 U980 ( .IN1(n913), .IN2(n955), .IN3(n929), .Q(n954) );
  INVX0 U981 ( .INP(n935), .ZN(n913) );
  OA21X1 U982 ( .IN1(n921), .IN2(n949), .IN3(n956), .Q(n923) );
  INVX0 U983 ( .INP(n930), .ZN(n949) );
  NAND2X0 U984 ( .IN1(n955), .IN2(n952), .QN(n930) );
  NAND2X0 U985 ( .IN1(keyinput121), .IN2(n918), .QN(n941) );
  MUX21X1 U986 ( .IN1(n957), .IN2(n958), .S(n959), .Q(n908) );
  NOR2X0 U987 ( .IN1(n960), .IN2(n961), .QN(n959) );
  AND3X1 U988 ( .IN1(N566), .IN2(n962), .IN3(n931), .Q(n960) );
  XOR3X1 U989 ( .IN1(keyinput127), .IN2(n963), .IN3(n964), .Q(n958) );
  XNOR2X1 U990 ( .IN1(n965), .IN2(n966), .Q(n964) );
  OA21X1 U991 ( .IN1(n967), .IN2(n968), .IN3(n969), .Q(n963) );
  XOR2X1 U992 ( .IN1(n970), .IN2(keyinput118), .Q(n969) );
  NAND2X0 U993 ( .IN1(n967), .IN2(n968), .QN(n970) );
  XNOR3X1 U994 ( .IN1(n971), .IN2(n972), .IN3(n973), .Q(n967) );
  NAND3X0 U995 ( .IN1(n974), .IN2(n975), .IN3(n976), .QN(n973) );
  XOR2X1 U996 ( .IN1(keyinput73), .IN2(n977), .Q(n976) );
  NOR2X0 U997 ( .IN1(n978), .IN2(n979), .QN(n977) );
  NAND3X0 U998 ( .IN1(N468), .IN2(n980), .IN3(n981), .QN(n974) );
  XOR3X1 U999 ( .IN1(n966), .IN2(n965), .IN3(n982), .Q(n957) );
  XOR3X1 U1000 ( .IN1(keyinput126), .IN2(keyinput122), .IN3(n983), .Q(n982) );
  OA21X1 U1001 ( .IN1(n968), .IN2(n984), .IN3(n985), .Q(n983) );
  XOR2X1 U1002 ( .IN1(keyinput117), .IN2(n986), .Q(n985) );
  AND2X1 U1003 ( .IN1(n968), .IN2(n984), .Q(n986) );
  XNOR3X1 U1004 ( .IN1(n987), .IN2(n988), .IN3(n989), .Q(n984) );
  XOR2X1 U1005 ( .IN1(n990), .IN2(n978), .Q(n965) );
  AO222X1 U1006 ( .IN1(n855), .IN2(n859), .IN3(N619), .IN4(n991), .IN5(N120), 
        .IN6(N625), .Q(N8075) );
  NAND2X0 U1007 ( .IN1(n858), .IN2(n907), .QN(n991) );
  XOR2X1 U1008 ( .IN1(n992), .IN2(n993), .Q(n858) );
  MUX21X1 U1009 ( .IN1(n994), .IN2(n995), .S(N583), .Q(n993) );
  XNOR3X1 U1010 ( .IN1(n996), .IN2(n997), .IN3(n998), .Q(n995) );
  XNOR3X1 U1011 ( .IN1(n999), .IN2(n1000), .IN3(n1001), .Q(n998) );
  AO22X1 U1012 ( .IN1(n1002), .IN2(n1003), .IN3(n1004), .IN4(n1005), .Q(n1001)
         );
  INVX0 U1013 ( .INP(n1006), .ZN(n1005) );
  OA21X1 U1014 ( .IN1(n1007), .IN2(n996), .IN3(n1008), .Q(n1004) );
  OA21X1 U1015 ( .IN1(n1009), .IN2(n1006), .IN3(n1010), .Q(n1002) );
  NOR2X0 U1016 ( .IN1(n1007), .IN2(n996), .QN(n1009) );
  OA21X1 U1017 ( .IN1(n1000), .IN2(n1010), .IN3(n1011), .Q(n999) );
  XNOR3X1 U1018 ( .IN1(n1006), .IN2(n997), .IN3(n1012), .Q(n994) );
  XNOR3X1 U1019 ( .IN1(n1003), .IN2(n1013), .IN3(n1011), .Q(n1012) );
  INVX0 U1020 ( .INP(n1014), .ZN(n997) );
  MUX21X1 U1021 ( .IN1(n1015), .IN2(n1016), .S(n1017), .Q(n1014) );
  OA21X1 U1022 ( .IN1(n1018), .IN2(n1019), .IN3(n1020), .Q(n1016) );
  XNOR2X1 U1023 ( .IN1(n1007), .IN2(n1021), .Q(n1015) );
  NAND2X0 U1024 ( .IN1(n1022), .IN2(n1023), .QN(n1006) );
  XNOR2X1 U1025 ( .IN1(n1024), .IN2(keyinput77), .Q(n1022) );
  MUX21X1 U1026 ( .IN1(n1025), .IN2(n1026), .S(n1027), .Q(n992) );
  AOI21X1 U1027 ( .IN1(N583), .IN2(n1028), .IN3(n1029), .QN(n1027) );
  XOR2X1 U1028 ( .IN1(keyinput85), .IN2(n1030), .Q(n1028) );
  AO21X1 U1029 ( .IN1(n1031), .IN2(n1032), .IN3(n1033), .Q(n1026) );
  XOR2X1 U1030 ( .IN1(keyinput124), .IN2(n1034), .Q(n1033) );
  NOR2X0 U1031 ( .IN1(n1032), .IN2(n1031), .QN(n1034) );
  XOR3X1 U1032 ( .IN1(n1035), .IN2(n1036), .IN3(n1037), .Q(n1031) );
  XNOR3X1 U1033 ( .IN1(n1038), .IN2(n1039), .IN3(n1040), .Q(n1037) );
  NOR2X0 U1034 ( .IN1(keyinput119), .IN2(n1041), .QN(n1038) );
  XOR2X1 U1035 ( .IN1(n1042), .IN2(n1043), .Q(n1035) );
  XNOR3X1 U1036 ( .IN1(n1040), .IN2(n1044), .IN3(n1045), .Q(n1025) );
  XNOR3X1 U1037 ( .IN1(n1046), .IN2(n1032), .IN3(n1047), .Q(n1045) );
  NAND2X0 U1038 ( .IN1(keyinput86), .IN2(n1048), .QN(n1047) );
  XOR2X1 U1039 ( .IN1(n1049), .IN2(n1050), .Q(n1048) );
  MUX21X1 U1040 ( .IN1(n1051), .IN2(n1042), .S(n1052), .Q(n1050) );
  NOR2X0 U1041 ( .IN1(n1053), .IN2(n1042), .QN(n1051) );
  AO21X1 U1042 ( .IN1(n1043), .IN2(n1054), .IN3(n1055), .Q(n1042) );
  NOR2X0 U1043 ( .IN1(n1056), .IN2(n1036), .QN(n1049) );
  NAND2X0 U1044 ( .IN1(n1057), .IN2(n1058), .QN(n1036) );
  XNOR3X1 U1045 ( .IN1(n1059), .IN2(n1060), .IN3(n1061), .Q(n859) );
  XNOR2X1 U1046 ( .IN1(keyinput83), .IN2(n1062), .Q(n1061) );
  OA21X1 U1047 ( .IN1(n1063), .IN2(n1064), .IN3(n1065), .Q(n1062) );
  XOR2X1 U1048 ( .IN1(n1066), .IN2(keyinput79), .Q(n1065) );
  NAND3X0 U1049 ( .IN1(n1067), .IN2(n1068), .IN3(n1064), .QN(n1066) );
  XNOR2X1 U1050 ( .IN1(n1069), .IN2(n1070), .Q(n1064) );
  NAND2X0 U1051 ( .IN1(n1071), .IN2(keyinput45), .QN(n1069) );
  MUX21X1 U1052 ( .IN1(n877), .IN2(n878), .S(n1072), .Q(n1071) );
  AND2X1 U1053 ( .IN1(n1068), .IN2(n1067), .Q(n1063) );
  NAND3X0 U1054 ( .IN1(n1073), .IN2(n1074), .IN3(n1075), .QN(n1067) );
  XNOR2X1 U1055 ( .IN1(keyinput28), .IN2(n1076), .Q(n1075) );
  NAND2X0 U1056 ( .IN1(n1077), .IN2(n1078), .QN(n1068) );
  INVX0 U1057 ( .INP(n1073), .ZN(n1078) );
  NAND2X0 U1058 ( .IN1(n1079), .IN2(n1080), .QN(n1073) );
  XOR2X1 U1059 ( .IN1(n1081), .IN2(keyinput41), .Q(n1079) );
  NAND2X0 U1060 ( .IN1(n1082), .IN2(n1083), .QN(n1081) );
  MUX21X1 U1061 ( .IN1(n1076), .IN2(n1084), .S(keyinput28), .Q(n1077) );
  XNOR3X1 U1062 ( .IN1(n1085), .IN2(n1086), .IN3(n1087), .Q(n1060) );
  MUX21X1 U1063 ( .IN1(n1088), .IN2(n1089), .S(n1090), .Q(n1087) );
  XNOR2X1 U1064 ( .IN1(N242), .IN2(n1091), .Q(n1089) );
  XNOR2X1 U1065 ( .IN1(n1091), .IN2(n877), .Q(n1088) );
  MUX21X1 U1066 ( .IN1(n1092), .IN2(n1093), .S(N503), .Q(n1091) );
  MUX21X1 U1067 ( .IN1(n877), .IN2(n878), .S(n1094), .Q(n1093) );
  MUX21X1 U1068 ( .IN1(n1095), .IN2(n1096), .S(keyinput20), .Q(n1092) );
  NAND2X0 U1069 ( .IN1(N254), .IN2(n1094), .QN(n1096) );
  MUX21X1 U1070 ( .IN1(N242), .IN2(N254), .S(n1094), .Q(n1095) );
  MUX41X1 U1071 ( .IN1(N251), .IN3(n888), .IN2(N248), .IN4(n887), .S0(n1097), 
        .S1(N341), .Q(n1085) );
  OA21X1 U1072 ( .IN1(N534), .IN2(n1098), .IN3(n1099), .Q(n1059) );
  XOR2X1 U1073 ( .IN1(keyinput27), .IN2(n1100), .Q(n1099) );
  NOR2X0 U1074 ( .IN1(n1101), .IN2(n1102), .QN(n1100) );
  MUX21X1 U1075 ( .IN1(n878), .IN2(n877), .S(N351), .Q(n1102) );
  MUX21X1 U1076 ( .IN1(N254), .IN2(N242), .S(N351), .Q(n1098) );
  AO221X1 U1077 ( .IN1(n1103), .IN2(n1104), .IN3(n1105), .IN4(n1106), .IN5(
        n1107), .Q(N7761) );
  AO22X1 U1078 ( .IN1(N191), .IN2(n1108), .IN3(N161), .IN4(n1109), .Q(n1107)
         );
  AO221X1 U1079 ( .IN1(n1103), .IN2(n1110), .IN3(n1105), .IN4(n1111), .IN5(
        n1112), .Q(N7760) );
  AO22X1 U1080 ( .IN1(N194), .IN2(n1108), .IN3(N164), .IN4(n1109), .Q(n1112)
         );
  AO221X1 U1081 ( .IN1(n1103), .IN2(n1113), .IN3(n1105), .IN4(n1114), .IN5(
        n1115), .Q(N7759) );
  AO22X1 U1082 ( .IN1(N197), .IN2(n1108), .IN3(N167), .IN4(n1109), .Q(n1115)
         );
  AO221X1 U1083 ( .IN1(n1103), .IN2(n1116), .IN3(n1105), .IN4(n1117), .IN5(
        n1118), .Q(N7758) );
  AO22X1 U1084 ( .IN1(N203), .IN2(n1108), .IN3(N173), .IN4(n1109), .Q(n1118)
         );
  AO221X1 U1085 ( .IN1(n1119), .IN2(n1106), .IN3(n1120), .IN4(N191), .IN5(
        n1121), .Q(N7757) );
  AO222X1 U1086 ( .IN1(n1122), .IN2(keyinput4), .IN3(n1123), .IN4(keyinput113), 
        .IN5(N137), .IN6(n1124), .Q(n1121) );
  AO22X1 U1087 ( .IN1(n1125), .IN2(n1126), .IN3(n1127), .IN4(n1128), .Q(n1124)
         );
  INVX0 U1088 ( .INP(keyinput113), .ZN(n1128) );
  NAND3X0 U1089 ( .IN1(n1104), .IN2(n839), .IN3(N571), .QN(n1127) );
  INVX0 U1090 ( .INP(keyinput4), .ZN(n1126) );
  NAND3X0 U1091 ( .IN1(N571), .IN2(N574), .IN3(N161), .QN(n1125) );
  AND2X1 U1092 ( .IN1(n1104), .IN2(n1129), .Q(n1123) );
  AND2X1 U1093 ( .IN1(N161), .IN2(n1130), .Q(n1122) );
  AO221X1 U1094 ( .IN1(n1129), .IN2(n1110), .IN3(n1119), .IN4(n1111), .IN5(
        n1131), .Q(N7756) );
  AO22X1 U1095 ( .IN1(n1120), .IN2(N194), .IN3(n1130), .IN4(N164), .Q(n1131)
         );
  AO221X1 U1096 ( .IN1(n1129), .IN2(n1113), .IN3(n1119), .IN4(n1114), .IN5(
        n1132), .Q(N7755) );
  AO22X1 U1097 ( .IN1(n1120), .IN2(N197), .IN3(n1130), .IN4(N167), .Q(n1132)
         );
  AO221X1 U1098 ( .IN1(n1129), .IN2(n1116), .IN3(n1119), .IN4(n1117), .IN5(
        n1133), .Q(N7754) );
  AO22X1 U1099 ( .IN1(n1120), .IN2(N203), .IN3(n1130), .IN4(N173), .Q(n1133)
         );
  AO221X1 U1100 ( .IN1(n843), .IN2(n1116), .IN3(n1134), .IN4(n1117), .IN5(
        n1135), .Q(N7742) );
  AO22X1 U1101 ( .IN1(N40), .IN2(n845), .IN3(N91), .IN4(n1136), .Q(n1135) );
  AO221X1 U1102 ( .IN1(n843), .IN2(n1113), .IN3(n1134), .IN4(n1114), .IN5(
        n1137), .Q(N7741) );
  AO22X1 U1103 ( .IN1(N103), .IN2(n845), .IN3(N100), .IN4(n1136), .Q(n1137) );
  XNOR2X1 U1104 ( .IN1(keyinput120), .IN2(n1138), .Q(N7740) );
  OA221X1 U1105 ( .IN1(n1139), .IN2(n1140), .IN3(N7705), .IN4(n1141), .IN5(
        n1142), .Q(n1138) );
  AOI22X1 U1106 ( .IN1(n1136), .IN2(N46), .IN3(n1111), .IN4(n1134), .QN(n1142)
         );
  INVX0 U1107 ( .INP(N49), .ZN(n1140) );
  AO221X1 U1108 ( .IN1(n848), .IN2(n1116), .IN3(n847), .IN4(n1117), .IN5(n1143), .Q(N7739) );
  AO21X1 U1109 ( .IN1(N91), .IN2(n851), .IN3(n1144), .Q(n1143) );
  XOR2X1 U1110 ( .IN1(n1145), .IN2(keyinput6), .Q(n1144) );
  NAND2X0 U1111 ( .IN1(N40), .IN2(n850), .QN(n1145) );
  AO221X1 U1112 ( .IN1(n848), .IN2(n1113), .IN3(N100), .IN4(n851), .IN5(n1146), 
        .Q(N7738) );
  AO21X1 U1113 ( .IN1(N103), .IN2(n850), .IN3(n1147), .Q(n1146) );
  XOR2X1 U1114 ( .IN1(keyinput115), .IN2(n1148), .Q(n1147) );
  NOR2X0 U1115 ( .IN1(N7701), .IN2(n1149), .QN(n1148) );
  AO221X1 U1116 ( .IN1(n848), .IN2(n1110), .IN3(n847), .IN4(n1111), .IN5(n1150), .Q(N7737) );
  AO22X1 U1117 ( .IN1(N49), .IN2(n850), .IN3(N46), .IN4(n851), .Q(n1150) );
  AO221X1 U1118 ( .IN1(n848), .IN2(n1104), .IN3(n847), .IN4(n1106), .IN5(n1151), .Q(N7736) );
  AO22X1 U1119 ( .IN1(N106), .IN2(n850), .IN3(N109), .IN4(n851), .Q(n1151) );
  AO221X1 U1120 ( .IN1(n1134), .IN2(n1106), .IN3(N109), .IN4(n1136), .IN5(
        n1152), .Q(N7735) );
  AO21X1 U1121 ( .IN1(N106), .IN2(n845), .IN3(n1153), .Q(n1152) );
  XOR2X1 U1122 ( .IN1(n1154), .IN2(keyinput114), .Q(n1153) );
  NAND2X0 U1123 ( .IN1(n843), .IN2(n1104), .QN(n1154) );
  INVX0 U1124 ( .INP(n1116), .ZN(N7707) );
  AO222X1 U1125 ( .IN1(n1155), .IN2(n855), .IN3(n1156), .IN4(n852), .IN5(N113), 
        .IN6(n1157), .Q(n1116) );
  INVX0 U1126 ( .INP(n1113), .ZN(N7706) );
  AO222X1 U1127 ( .IN1(n1158), .IN2(n855), .IN3(n1159), .IN4(n852), .IN5(N53), 
        .IN6(n1157), .Q(n1113) );
  INVX0 U1128 ( .INP(n1110), .ZN(N7705) );
  AO222X1 U1129 ( .IN1(n1160), .IN2(n855), .IN3(n852), .IN4(n1161), .IN5(N114), 
        .IN6(n1157), .Q(n1110) );
  XNOR2X1 U1130 ( .IN1(keyinput116), .IN2(n1104), .Q(N7704) );
  AO221X1 U1131 ( .IN1(n852), .IN2(n1162), .IN3(n855), .IN4(n902), .IN5(n1163), 
        .Q(n1104) );
  XNOR2X1 U1132 ( .IN1(n1164), .IN2(keyinput33), .Q(n1163) );
  NAND2X0 U1133 ( .IN1(N115), .IN2(n1157), .QN(n1164) );
  NOR4X0 U1134 ( .IN1(n1165), .IN2(N1152), .IN3(N1155), .IN4(N1153), .QN(N7703) );
  NAND3X0 U1135 ( .IN1(N556), .IN2(N386), .IN3(n1166), .QN(n1165) );
  XOR2X1 U1136 ( .IN1(n1167), .IN2(keyinput111), .Q(n1166) );
  OR4X1 U1137 ( .IN1(N7474), .IN2(N7476), .IN3(N6716), .IN4(n1168), .Q(n1167)
         );
  OR2X1 U1138 ( .IN1(N6877), .IN2(n1169), .Q(n1168) );
  INVX0 U1139 ( .INP(n1117), .ZN(N7702) );
  AO222X1 U1140 ( .IN1(n1170), .IN2(n852), .IN3(n1171), .IN4(n855), .IN5(N112), 
        .IN6(n1157), .Q(n1117) );
  INVX0 U1141 ( .INP(n1114), .ZN(N7701) );
  AO222X1 U1142 ( .IN1(n1172), .IN2(n855), .IN3(n852), .IN4(n1173), .IN5(N116), 
        .IN6(n1157), .Q(n1114) );
  INVX0 U1143 ( .INP(n1111), .ZN(N7700) );
  AO222X1 U1144 ( .IN1(n855), .IN2(n1174), .IN3(n852), .IN4(n1175), .IN5(N121), 
        .IN6(n1157), .Q(n1111) );
  INVX0 U1145 ( .INP(n1106), .ZN(N7699) );
  AO222X1 U1146 ( .IN1(n855), .IN2(n1176), .IN3(n852), .IN4(n1177), .IN5(N123), 
        .IN6(n1157), .Q(n1106) );
  XNOR2X1 U1147 ( .IN1(N7432), .IN2(n1178), .Q(N7698) );
  AOI21X1 U1148 ( .IN1(N631), .IN2(N135), .IN3(n1179), .QN(N7626) );
  INVX0 U1149 ( .INP(n1180), .ZN(n1179) );
  MUX41X1 U1150 ( .IN1(n1176), .IN3(n1178), .IN2(N123), .IN4(n1177), .S0(N603), 
        .S1(N599), .Q(n1180) );
  XOR2X1 U1151 ( .IN1(n1044), .IN2(N132), .Q(n1178) );
  AO221X1 U1152 ( .IN1(N149), .IN2(n1108), .IN3(n1105), .IN4(n1181), .IN5(
        n1182), .Q(N7607) );
  AO22X1 U1153 ( .IN1(N146), .IN2(n1109), .IN3(n1103), .IN4(n1183), .Q(n1182)
         );
  AO221X1 U1154 ( .IN1(N155), .IN2(n1108), .IN3(n1105), .IN4(n1184), .IN5(
        n1185), .Q(N7606) );
  AO22X1 U1155 ( .IN1(N152), .IN2(n1109), .IN3(n1103), .IN4(n1186), .Q(n1185)
         );
  AO221X1 U1156 ( .IN1(n1103), .IN2(n1187), .IN3(N188), .IN4(n1108), .IN5(
        n1188), .Q(N7605) );
  AO21X1 U1157 ( .IN1(n1105), .IN2(n1189), .IN3(n1190), .Q(n1188) );
  MUX21X1 U1158 ( .IN1(n1191), .IN2(n1192), .S(keyinput5), .Q(n1190) );
  NOR2X0 U1159 ( .IN1(n1193), .IN2(n1194), .QN(n1192) );
  AND3X1 U1160 ( .IN1(N580), .IN2(N577), .IN3(N158), .Q(n1193) );
  AND2X1 U1161 ( .IN1(n1109), .IN2(N158), .Q(n1191) );
  AO221X1 U1162 ( .IN1(n1103), .IN2(n1195), .IN3(N170), .IN4(n1109), .IN5(
        n1196), .Q(N7604) );
  AO21X1 U1163 ( .IN1(n1108), .IN2(N200), .IN3(n1197), .Q(n1196) );
  INVX0 U1164 ( .INP(n1198), .ZN(n1197) );
  MUX21X1 U1165 ( .IN1(n1199), .IN2(n1200), .S(keyinput107), .Q(n1198) );
  NAND2X0 U1166 ( .IN1(n1105), .IN2(n1201), .QN(n1200) );
  NAND2X0 U1167 ( .IN1(N137), .IN2(n1202), .QN(n1199) );
  OR3X1 U1168 ( .IN1(N577), .IN2(N580), .IN3(N7465), .Q(n1202) );
  AO221X1 U1169 ( .IN1(N149), .IN2(n1120), .IN3(n1119), .IN4(n1181), .IN5(
        n1203), .Q(N7603) );
  AO22X1 U1170 ( .IN1(N146), .IN2(n1130), .IN3(n1129), .IN4(n1183), .Q(n1203)
         );
  AO221X1 U1171 ( .IN1(N155), .IN2(n1120), .IN3(n1119), .IN4(n1184), .IN5(
        n1204), .Q(N7602) );
  AO22X1 U1172 ( .IN1(N152), .IN2(n1130), .IN3(n1129), .IN4(n1186), .Q(n1204)
         );
  AO221X1 U1173 ( .IN1(n1129), .IN2(n1187), .IN3(N158), .IN4(n1130), .IN5(
        n1205), .Q(N7601) );
  AO22X1 U1174 ( .IN1(n1119), .IN2(n1189), .IN3(N188), .IN4(n1120), .Q(n1205)
         );
  AO221X1 U1175 ( .IN1(n1129), .IN2(n1195), .IN3(N170), .IN4(n1130), .IN5(
        n1206), .Q(N7600) );
  AO22X1 U1176 ( .IN1(n1119), .IN2(n1201), .IN3(N200), .IN4(n1120), .Q(n1206)
         );
  AO221X1 U1177 ( .IN1(n843), .IN2(n1187), .IN3(n842), .IN4(n1189), .IN5(n1207), .Q(N7522) );
  AO22X1 U1178 ( .IN1(N70), .IN2(n845), .IN3(N67), .IN4(n846), .Q(n1207) );
  AO221X1 U1179 ( .IN1(n842), .IN2(n1184), .IN3(N73), .IN4(n846), .IN5(n1208), 
        .Q(N7521) );
  AO21X1 U1180 ( .IN1(N17), .IN2(n845), .IN3(n1209), .Q(n1208) );
  XOR2X1 U1181 ( .IN1(keyinput109), .IN2(n1210), .Q(n1209) );
  NOR2X0 U1182 ( .IN1(N7472), .IN2(n1141), .QN(n1210) );
  INVX0 U1183 ( .INP(n843), .ZN(n1141) );
  AO221X1 U1184 ( .IN1(n843), .IN2(n1183), .IN3(n842), .IN4(n1181), .IN5(n1211), .Q(N7520) );
  AO22X1 U1185 ( .IN1(N20), .IN2(n845), .IN3(N76), .IN4(n846), .Q(n1211) );
  AO221X1 U1186 ( .IN1(N43), .IN2(n1136), .IN3(n843), .IN4(n1195), .IN5(n1212), 
        .Q(N7519) );
  AO21X1 U1187 ( .IN1(N37), .IN2(n845), .IN3(n1213), .Q(n1212) );
  XOR2X1 U1188 ( .IN1(n1214), .IN2(keyinput108), .Q(n1213) );
  NAND2X0 U1189 ( .IN1(n1134), .IN2(n1201), .QN(n1214) );
  AO221X1 U1190 ( .IN1(n848), .IN2(n1187), .IN3(N67), .IN4(n851), .IN5(n1215), 
        .Q(N7518) );
  AO21X1 U1191 ( .IN1(N70), .IN2(n850), .IN3(n1216), .Q(n1215) );
  XOR2X1 U1192 ( .IN1(keyinput103), .IN2(n1217), .Q(n1216) );
  NOR2X0 U1193 ( .IN1(N7363), .IN2(n1149), .QN(n1217) );
  INVX0 U1194 ( .INP(n847), .ZN(n1149) );
  AO221X1 U1195 ( .IN1(n848), .IN2(n1186), .IN3(n847), .IN4(n1184), .IN5(n1218), .Q(N7517) );
  AO22X1 U1196 ( .IN1(N17), .IN2(n850), .IN3(N73), .IN4(n851), .Q(n1218) );
  AO221X1 U1197 ( .IN1(n848), .IN2(n1183), .IN3(n847), .IN4(n1181), .IN5(n1219), .Q(N7516) );
  AO22X1 U1198 ( .IN1(N20), .IN2(n850), .IN3(N76), .IN4(n851), .Q(n1219) );
  AO221X1 U1199 ( .IN1(N182), .IN2(n1108), .IN3(n1105), .IN4(n1220), .IN5(
        n1221), .Q(N7511) );
  AO22X1 U1200 ( .IN1(N185), .IN2(n1109), .IN3(n1103), .IN4(n1222), .Q(n1221)
         );
  NOR3X0 U1201 ( .IN1(n831), .IN2(N580), .IN3(n1194), .QN(n1103) );
  AND3X1 U1202 ( .IN1(N580), .IN2(N577), .IN3(N137), .Q(n1109) );
  NOR3X0 U1203 ( .IN1(N577), .IN2(N580), .IN3(n1194), .QN(n1105) );
  AND3X1 U1204 ( .IN1(N580), .IN2(n831), .IN3(N137), .Q(n1108) );
  INVX0 U1205 ( .INP(N577), .ZN(n831) );
  AO221X1 U1206 ( .IN1(N182), .IN2(n1120), .IN3(n1119), .IN4(n1220), .IN5(
        n1223), .Q(N7506) );
  AO22X1 U1207 ( .IN1(N185), .IN2(n1130), .IN3(n1129), .IN4(n1222), .Q(n1223)
         );
  AND3X1 U1208 ( .IN1(N137), .IN2(n839), .IN3(N571), .Q(n1129) );
  NOR3X0 U1209 ( .IN1(n839), .IN2(n1194), .IN3(n840), .QN(n1130) );
  AND3X1 U1210 ( .IN1(n840), .IN2(n839), .IN3(N137), .Q(n1119) );
  INVX0 U1211 ( .INP(N571), .ZN(n840) );
  NOR2X0 U1212 ( .IN1(n835), .IN2(n1194), .QN(n1120) );
  INVX0 U1213 ( .INP(N137), .ZN(n1194) );
  INVX0 U1214 ( .INP(n841), .ZN(n835) );
  NOR2X0 U1215 ( .IN1(n839), .IN2(N571), .QN(n841) );
  INVX0 U1216 ( .INP(N574), .ZN(n839) );
  NOR4X0 U1217 ( .IN1(n1224), .IN2(n1225), .IN3(n1177), .IN4(n1175), .QN(N7504) );
  INVX0 U1218 ( .INP(n1226), .ZN(n1175) );
  MUX21X1 U1219 ( .IN1(n1227), .IN2(n1228), .S(n1229), .Q(n1226) );
  OA21X1 U1220 ( .IN1(n1230), .IN2(n1231), .IN3(n1232), .Q(n1228) );
  OA21X1 U1221 ( .IN1(keyinput88), .IN2(n1233), .IN3(n1234), .Q(n1227) );
  AO22X1 U1222 ( .IN1(n1230), .IN2(n1235), .IN3(n1231), .IN4(n1236), .Q(n1234)
         );
  INVX0 U1223 ( .INP(keyinput88), .ZN(n1236) );
  INVX0 U1224 ( .INP(N7432), .ZN(n1177) );
  OR3X1 U1225 ( .IN1(n1237), .IN2(n1170), .IN3(n1238), .Q(n1225) );
  XNOR2X1 U1226 ( .IN1(n1046), .IN2(n1229), .Q(n1170) );
  NAND4X0 U1227 ( .IN1(n1239), .IN2(n1240), .IN3(n1241), .IN4(n1242), .QN(
        n1224) );
  INVX0 U1228 ( .INP(n1243), .ZN(n1242) );
  XNOR2X1 U1229 ( .IN1(n1244), .IN2(keyinput97), .Q(n1241) );
  XNOR2X1 U1230 ( .IN1(n1173), .IN2(keyinput106), .Q(n1240) );
  INVX0 U1231 ( .INP(n1245), .ZN(n1173) );
  MUX21X1 U1232 ( .IN1(n1246), .IN2(n1247), .S(n1229), .Q(n1245) );
  OA21X1 U1233 ( .IN1(n1043), .IN2(n1248), .IN3(n1249), .Q(n1247) );
  XOR2X1 U1234 ( .IN1(n1250), .IN2(keyinput89), .Q(n1249) );
  NAND2X0 U1235 ( .IN1(n1043), .IN2(n1248), .QN(n1250) );
  XNOR3X1 U1236 ( .IN1(keyinput93), .IN2(n1251), .IN3(n1252), .Q(n1246) );
  NAND2X0 U1237 ( .IN1(keyinput84), .IN2(n1052), .QN(n1252) );
  XNOR2X1 U1238 ( .IN1(n1253), .IN2(keyinput98), .Q(n1239) );
  NOR4X0 U1239 ( .IN1(n1254), .IN2(n1255), .IN3(n1256), .IN4(n1257), .QN(N7503) );
  OR3X1 U1240 ( .IN1(n1156), .IN2(n1159), .IN3(n1258), .Q(n1255) );
  AND2X1 U1241 ( .IN1(n1259), .IN2(n979), .Q(n1159) );
  MUX21X1 U1242 ( .IN1(n1260), .IN2(n1261), .S(n966), .Q(n1259) );
  NAND2X0 U1243 ( .IN1(n1262), .IN2(n1263), .QN(n1261) );
  OA21X1 U1244 ( .IN1(n971), .IN2(n1263), .IN3(n1262), .Q(n1260) );
  INVX0 U1245 ( .INP(n987), .ZN(n1262) );
  XNOR2X1 U1246 ( .IN1(n1263), .IN2(n968), .Q(n1156) );
  INVX0 U1247 ( .INP(n1264), .ZN(n968) );
  OR4X1 U1248 ( .IN1(n1161), .IN2(n1162), .IN3(n1265), .IN4(n1266), .Q(n1254)
         );
  XOR2X1 U1249 ( .IN1(n1267), .IN2(n1268), .Q(n1162) );
  OA21X1 U1250 ( .IN1(n1269), .IN2(n989), .IN3(n1270), .Q(n1268) );
  NOR2X0 U1251 ( .IN1(n1271), .IN2(n1272), .QN(n989) );
  INVX0 U1252 ( .INP(n1263), .ZN(n1269) );
  INVX0 U1253 ( .INP(n1273), .ZN(n1161) );
  MUX21X1 U1254 ( .IN1(n1274), .IN2(n1275), .S(n1263), .Q(n1273) );
  AO21X1 U1255 ( .IN1(N4), .IN2(n1276), .IN3(n1277), .Q(n1263) );
  XNOR2X1 U1256 ( .IN1(n988), .IN2(n981), .Q(n1275) );
  NAND2X0 U1257 ( .IN1(n972), .IN2(n1278), .QN(n988) );
  AO21X1 U1258 ( .IN1(n972), .IN2(n978), .IN3(n1279), .Q(n1274) );
  XOR2X1 U1259 ( .IN1(n1280), .IN2(keyinput92), .Q(n1279) );
  NAND2X0 U1260 ( .IN1(n981), .IN2(n1281), .QN(n1280) );
  AO21X1 U1261 ( .IN1(n1282), .IN2(n1283), .IN3(n1284), .Q(N7476) );
  XOR2X1 U1262 ( .IN1(n1285), .IN2(keyinput99), .Q(n1284) );
  OR2X1 U1263 ( .IN1(n1283), .IN2(n1282), .Q(n1285) );
  NAND2X0 U1264 ( .IN1(n1286), .IN2(n1287), .QN(n1283) );
  NAND3X0 U1265 ( .IN1(n1288), .IN2(n1289), .IN3(n1290), .QN(n1287) );
  XNOR2X1 U1266 ( .IN1(keyinput82), .IN2(n1291), .Q(n1286) );
  AOI21X1 U1267 ( .IN1(n1288), .IN2(n1290), .IN3(n1289), .QN(n1291) );
  AO21X1 U1268 ( .IN1(n1292), .IN2(n1293), .IN3(n1294), .Q(n1289) );
  XOR2X1 U1269 ( .IN1(n1295), .IN2(keyinput65), .Q(n1294) );
  OR2X1 U1270 ( .IN1(n1293), .IN2(n1292), .Q(n1295) );
  XOR2X1 U1271 ( .IN1(n1296), .IN2(keyinput64), .Q(n1290) );
  NAND2X0 U1272 ( .IN1(n1297), .IN2(n932), .QN(n1296) );
  OR2X1 U1273 ( .IN1(n932), .IN2(n1297), .Q(n1288) );
  INVX0 U1274 ( .INP(n1298), .ZN(n1297) );
  XOR2X1 U1275 ( .IN1(n1299), .IN2(n1300), .Q(n1282) );
  XOR3X1 U1276 ( .IN1(n1301), .IN2(n1302), .IN3(n1303), .Q(n1300) );
  XOR2X1 U1277 ( .IN1(n1304), .IN2(n980), .Q(n1303) );
  XOR3X1 U1278 ( .IN1(keyinput95), .IN2(keyinput71), .IN3(n1305), .Q(n1299) );
  XOR2X1 U1279 ( .IN1(n1306), .IN2(n1307), .Q(n1305) );
  AO22X1 U1280 ( .IN1(N292), .IN2(N335), .IN3(N289), .IN4(n1308), .Q(n1306) );
  AO21X1 U1281 ( .IN1(n1309), .IN2(n1310), .IN3(n1311), .Q(N7474) );
  XOR2X1 U1282 ( .IN1(keyinput102), .IN2(n1312), .Q(n1311) );
  NOR2X0 U1283 ( .IN1(n1309), .IN2(n1310), .QN(n1312) );
  XNOR3X1 U1284 ( .IN1(n1313), .IN2(n1314), .IN3(n1315), .Q(n1310) );
  XNOR2X1 U1285 ( .IN1(n1044), .IN2(n1316), .Q(n1315) );
  XNOR3X1 U1286 ( .IN1(n1317), .IN2(n1318), .IN3(n1319), .Q(n1309) );
  AO22X1 U1287 ( .IN1(N372), .IN2(N332), .IN3(N369), .IN4(n1320), .Q(n1319) );
  NOR2X0 U1288 ( .IN1(keyinput78), .IN2(n1321), .QN(n1318) );
  XNOR3X1 U1289 ( .IN1(n1322), .IN2(n1323), .IN3(n1324), .Q(n1321) );
  NAND2X0 U1290 ( .IN1(keyinput59), .IN2(n1325), .QN(n1324) );
  OA21X1 U1291 ( .IN1(n1326), .IN2(n1327), .IN3(n1328), .Q(n1323) );
  XOR2X1 U1292 ( .IN1(n1329), .IN2(keyinput60), .Q(n1328) );
  NAND2X0 U1293 ( .IN1(n1327), .IN2(n1326), .QN(n1329) );
  INVX0 U1294 ( .INP(n1187), .ZN(N7473) );
  AO222X1 U1295 ( .IN1(n1330), .IN2(n855), .IN3(n1256), .IN4(n852), .IN5(N126), 
        .IN6(n1157), .Q(n1187) );
  XOR2X1 U1296 ( .IN1(n1331), .IN2(n933), .Q(n1256) );
  INVX0 U1297 ( .INP(n1186), .ZN(N7472) );
  AO222X1 U1298 ( .IN1(n1332), .IN2(n855), .IN3(n852), .IN4(n1266), .IN5(N127), 
        .IN6(n1157), .Q(n1186) );
  XOR2X1 U1299 ( .IN1(n1333), .IN2(n1334), .Q(n1266) );
  INVX0 U1300 ( .INP(n1183), .ZN(N7471) );
  AO222X1 U1301 ( .IN1(n1335), .IN2(n855), .IN3(n1258), .IN4(n852), .IN5(N128), 
        .IN6(n1157), .Q(n1183) );
  XOR2X1 U1302 ( .IN1(n1336), .IN2(n917), .Q(n1258) );
  INVX0 U1303 ( .INP(n1195), .ZN(N7470) );
  AO221X1 U1304 ( .IN1(n842), .IN2(n1220), .IN3(N11), .IN4(n846), .IN5(n1337), 
        .Q(N7469) );
  AO22X1 U1305 ( .IN1(N61), .IN2(n845), .IN3(n843), .IN4(n1222), .Q(n1337) );
  MUX21X1 U1306 ( .IN1(n845), .IN2(n1136), .S(keyinput7), .Q(n846) );
  AND2X1 U1307 ( .IN1(N616), .IN2(n1338), .Q(n1136) );
  INVX0 U1308 ( .INP(n1139), .ZN(n845) );
  NAND2X0 U1309 ( .IN1(N616), .IN2(N613), .QN(n1139) );
  MUX21X1 U1310 ( .IN1(n843), .IN2(n1134), .S(keyinput7), .Q(n842) );
  NOR2X0 U1311 ( .IN1(N613), .IN2(N616), .QN(n1134) );
  NOR2X0 U1312 ( .IN1(n1338), .IN2(N616), .QN(n843) );
  INVX0 U1313 ( .INP(N613), .ZN(n1338) );
  INVX0 U1314 ( .INP(n1184), .ZN(N7467) );
  AO221X1 U1315 ( .IN1(n1339), .IN2(n855), .IN3(N119), .IN4(n1157), .IN5(n1340), .Q(n1184) );
  XOR2X1 U1316 ( .IN1(n1341), .IN2(keyinput100), .Q(n1340) );
  NAND2X0 U1317 ( .IN1(n852), .IN2(n1244), .QN(n1341) );
  XNOR2X1 U1318 ( .IN1(n1342), .IN2(n1019), .Q(n1244) );
  INVX0 U1319 ( .INP(n1181), .ZN(N7466) );
  AO221X1 U1320 ( .IN1(n1237), .IN2(n852), .IN3(N130), .IN4(n1157), .IN5(n1343), .Q(n1181) );
  XOR2X1 U1321 ( .IN1(keyinput42), .IN2(n1344), .Q(n1343) );
  AND2X1 U1322 ( .IN1(n1345), .IN2(n855), .Q(n1344) );
  XNOR2X1 U1323 ( .IN1(n1346), .IN2(n1347), .Q(n1237) );
  NAND2X0 U1324 ( .IN1(keyinput90), .IN2(n1348), .QN(n1347) );
  NAND4X0 U1325 ( .IN1(n1349), .IN2(n1350), .IN3(n1351), .IN4(n1352), .QN(
        n1346) );
  NAND2X0 U1326 ( .IN1(N54), .IN2(n1353), .QN(n1350) );
  XNOR2X1 U1327 ( .IN1(keyinput76), .IN2(n1354), .Q(n1349) );
  INVX0 U1328 ( .INP(n1201), .ZN(N7465) );
  AO221X1 U1329 ( .IN1(n848), .IN2(n1222), .IN3(n847), .IN4(n1220), .IN5(n1355), .Q(N7449) );
  AO22X1 U1330 ( .IN1(N61), .IN2(n850), .IN3(N11), .IN4(n851), .Q(n1355) );
  MUX21X1 U1331 ( .IN1(n1356), .IN2(n1357), .S(n1229), .Q(N7432) );
  AND2X1 U1332 ( .IN1(n1358), .IN2(n1359), .Q(n1229) );
  NAND4X0 U1333 ( .IN1(N54), .IN2(n1360), .IN3(n1017), .IN4(n1348), .QN(n1359)
         );
  XNOR2X1 U1334 ( .IN1(n1232), .IN2(n1044), .Q(n1357) );
  XNOR2X1 U1335 ( .IN1(n1233), .IN2(n1044), .Q(n1356) );
  NAND2X0 U1336 ( .IN1(n1361), .IN2(n1235), .QN(n1233) );
  XNOR2X1 U1337 ( .IN1(keyinput104), .IN2(n1222), .Q(N7365) );
  AO221X1 U1338 ( .IN1(n852), .IN2(n1265), .IN3(N117), .IN4(n1157), .IN5(n1362), .Q(n1222) );
  XOR2X1 U1339 ( .IN1(n1363), .IN2(keyinput54), .Q(n1362) );
  NAND2X0 U1340 ( .IN1(n1364), .IN2(n855), .QN(n1363) );
  XOR2X1 U1341 ( .IN1(N4), .IN2(n918), .Q(n1265) );
  INVX0 U1342 ( .INP(n1189), .ZN(N7363) );
  AO222X1 U1343 ( .IN1(n1365), .IN2(n855), .IN3(n1238), .IN4(n852), .IN5(N129), 
        .IN6(n1157), .Q(n1189) );
  XNOR2X1 U1344 ( .IN1(n1366), .IN2(n1018), .Q(n1238) );
  INVX0 U1345 ( .INP(n1220), .ZN(N7015) );
  AO222X1 U1346 ( .IN1(n855), .IN2(n1086), .IN3(n852), .IN4(n1243), .IN5(N131), 
        .IN6(n1157), .Q(n1220) );
  AO21X1 U1347 ( .IN1(N54), .IN2(n996), .IN3(n1366), .Q(n1243) );
  NAND4X0 U1348 ( .IN1(n1057), .IN2(n1367), .IN3(n1044), .IN4(n1368), .QN(
        N6927) );
  NAND2X0 U1349 ( .IN1(n1056), .IN2(n1029), .QN(n1368) );
  XOR2X1 U1350 ( .IN1(keyinput81), .IN2(n1369), .Q(n1029) );
  OA21X1 U1351 ( .IN1(n1011), .IN2(n1370), .IN3(n1371), .Q(n1369) );
  OA221X1 U1352 ( .IN1(n1000), .IN2(n1352), .IN3(n1372), .IN4(n1000), .IN5(
        n1373), .Q(n1011) );
  AND2X1 U1353 ( .IN1(n1351), .IN2(n1354), .Q(n1372) );
  INVX0 U1354 ( .INP(n1013), .ZN(n1000) );
  INVX0 U1355 ( .INP(n1374), .ZN(n1056) );
  XNOR2X1 U1356 ( .IN1(keyinput72), .IN2(n1058), .Q(n1367) );
  NAND3X0 U1357 ( .IN1(n1032), .IN2(n1054), .IN3(n1043), .QN(n1058) );
  AOI21X1 U1358 ( .IN1(n1055), .IN2(n1032), .IN3(n1313), .QN(n1057) );
  AO21X1 U1359 ( .IN1(n1375), .IN2(n1376), .IN3(n1377), .Q(N6926) );
  AO21X1 U1360 ( .IN1(n1272), .IN2(n1277), .IN3(n1271), .Q(n1376) );
  AO21X1 U1361 ( .IN1(n1378), .IN2(n1379), .IN3(n1380), .Q(n1277) );
  NAND2X0 U1362 ( .IN1(n956), .IN2(n1381), .QN(n1379) );
  NAND3X0 U1363 ( .IN1(n940), .IN2(n1382), .IN3(n1334), .QN(n1381) );
  NAND2X0 U1364 ( .IN1(n952), .IN2(n1383), .QN(n1382) );
  OA21X1 U1365 ( .IN1(n929), .IN2(n917), .IN3(n1384), .Q(n956) );
  NAND3X0 U1366 ( .IN1(n1044), .IN2(n1385), .IN3(n1361), .QN(N6925) );
  INVX0 U1367 ( .INP(n1232), .ZN(n1361) );
  NAND2X0 U1368 ( .IN1(n1230), .IN2(n1231), .QN(n1232) );
  INVX0 U1369 ( .INP(n1313), .ZN(n1231) );
  AOI21X1 U1370 ( .IN1(n1043), .IN2(n1251), .IN3(n1055), .QN(n1230) );
  OR2X1 U1371 ( .IN1(n1235), .IN2(n1358), .Q(n1385) );
  OA21X1 U1372 ( .IN1(n1370), .IN2(n1386), .IN3(n1371), .Q(n1358) );
  NAND2X0 U1373 ( .IN1(N503), .IN2(n1327), .QN(n1371) );
  OA21X1 U1374 ( .IN1(n1387), .IN2(n1003), .IN3(n1373), .Q(n1386) );
  INVX0 U1375 ( .INP(n1008), .ZN(n1003) );
  NAND3X0 U1376 ( .IN1(n1351), .IN2(n1352), .IN3(n1354), .QN(n1008) );
  OR2X1 U1377 ( .IN1(n1023), .IN2(n1021), .Q(n1354) );
  NAND2X0 U1378 ( .IN1(n1024), .IN2(n1019), .QN(n1352) );
  NOR2X0 U1379 ( .IN1(n1007), .IN2(n1317), .QN(n1024) );
  INVX0 U1380 ( .INP(n996), .ZN(n1317) );
  NAND3X0 U1381 ( .IN1(n1388), .IN2(n1389), .IN3(n1390), .QN(N6924) );
  XNOR2X1 U1382 ( .IN1(n1391), .IN2(keyinput87), .Q(n1390) );
  NAND3X0 U1383 ( .IN1(n990), .IN2(n961), .IN3(n1272), .QN(n1391) );
  XOR2X1 U1384 ( .IN1(keyinput80), .IN2(n1392), .Q(n961) );
  OA221X1 U1385 ( .IN1(keyinput74), .IN2(n1393), .IN3(keyinput75), .IN4(n1394), 
        .IN5(n1395), .Q(n1392) );
  OA21X1 U1386 ( .IN1(n1396), .IN2(n912), .IN3(n1397), .Q(n1395) );
  XOR2X1 U1387 ( .IN1(keyinput49), .IN2(n1380), .Q(n1397) );
  AND2X1 U1388 ( .IN1(N435), .IN2(n1302), .Q(n1380) );
  OA221X1 U1389 ( .IN1(n1398), .IN2(n921), .IN3(n1399), .IN4(n1400), .IN5(
        n1384), .Q(n1396) );
  NAND2X0 U1390 ( .IN1(n1401), .IN2(n940), .QN(n1400) );
  INVX0 U1391 ( .INP(keyinput74), .ZN(n1399) );
  OA21X1 U1392 ( .IN1(n952), .IN2(n1402), .IN3(n955), .Q(n1398) );
  XNOR2X1 U1393 ( .IN1(n1383), .IN2(keyinput50), .Q(n955) );
  INVX0 U1394 ( .INP(keyinput75), .ZN(n1402) );
  NOR2X0 U1395 ( .IN1(n1403), .IN2(n952), .QN(n1394) );
  NAND2X0 U1396 ( .IN1(n953), .IN2(n933), .QN(n952) );
  INVX0 U1397 ( .INP(n962), .ZN(n1403) );
  NOR3X0 U1398 ( .IN1(n929), .IN2(n917), .IN3(n912), .QN(n1393) );
  INVX0 U1399 ( .INP(n1401), .ZN(n929) );
  INVX0 U1400 ( .INP(n1377), .ZN(n1389) );
  NAND2X0 U1401 ( .IN1(n990), .IN2(n1271), .QN(n1388) );
  INVX0 U1402 ( .INP(n1270), .ZN(n1271) );
  OA21X1 U1403 ( .IN1(n978), .IN2(n972), .IN3(n975), .Q(n1270) );
  INVX0 U1404 ( .INP(n1281), .ZN(n972) );
  AO21X1 U1405 ( .IN1(N468), .IN2(n980), .IN3(n1404), .Q(n1281) );
  INVX0 U1406 ( .INP(n979), .ZN(n1404) );
  NAND2X0 U1407 ( .IN1(n971), .IN2(n966), .QN(n979) );
  XOR3X1 U1408 ( .IN1(keyinput66), .IN2(n1405), .IN3(n1406), .Q(N6877) );
  AO221X1 U1409 ( .IN1(n1407), .IN2(n1408), .IN3(keyinput61), .IN4(n1409), 
        .IN5(n1410), .Q(n1406) );
  MUX21X1 U1410 ( .IN1(n1411), .IN2(n1412), .S(n1413), .Q(n1410) );
  OA21X1 U1411 ( .IN1(N265), .IN2(n886), .IN3(n1414), .Q(n1413) );
  XOR2X1 U1412 ( .IN1(keyinput22), .IN2(n1415), .Q(n1414) );
  NOR2X0 U1413 ( .IN1(N273), .IN2(n879), .QN(n1415) );
  INVX0 U1414 ( .INP(N273), .ZN(n886) );
  OAI22X1 U1415 ( .IN1(n1409), .IN2(keyinput61), .IN3(n1408), .IN4(n1407), 
        .QN(n1412) );
  NAND3X0 U1416 ( .IN1(n1416), .IN2(n1417), .IN3(keyinput55), .QN(n1411) );
  INVX0 U1417 ( .INP(keyinput61), .ZN(n1417) );
  XNOR2X1 U1418 ( .IN1(n1418), .IN2(n1419), .Q(n1416) );
  NAND2X0 U1419 ( .IN1(n1418), .IN2(n1419), .QN(n1409) );
  INVX0 U1420 ( .INP(keyinput55), .ZN(n1408) );
  OR2X1 U1421 ( .IN1(n1419), .IN2(n1418), .Q(n1407) );
  XOR2X1 U1422 ( .IN1(n1420), .IN2(N257), .Q(n1418) );
  NAND2X0 U1423 ( .IN1(keyinput16), .IN2(N234), .QN(n1420) );
  XOR3X1 U1424 ( .IN1(keyinput32), .IN2(n1421), .IN3(N289), .Q(n1419) );
  NOR2X0 U1425 ( .IN1(keyinput15), .IN2(n889), .QN(n1421) );
  INVX0 U1426 ( .INP(N281), .ZN(n889) );
  NOR2X0 U1427 ( .IN1(n1422), .IN2(n1423), .QN(n1405) );
  XOR2X1 U1428 ( .IN1(keyinput62), .IN2(n1424), .Q(n1423) );
  NOR2X0 U1429 ( .IN1(n1425), .IN2(n1426), .QN(n1424) );
  XNOR2X1 U1430 ( .IN1(N210), .IN2(n1427), .Q(n1426) );
  INVX0 U1431 ( .INP(n1428), .ZN(n1425) );
  XOR2X1 U1432 ( .IN1(keyinput56), .IN2(n1429), .Q(n1422) );
  NOR2X0 U1433 ( .IN1(n1430), .IN2(n1428), .QN(n1429) );
  XOR2X1 U1434 ( .IN1(N218), .IN2(N226), .Q(n1428) );
  XNOR2X1 U1435 ( .IN1(N206), .IN2(N210), .Q(n1430) );
  XNOR3X1 U1436 ( .IN1(n1431), .IN2(n1432), .IN3(n1433), .Q(N6716) );
  MUX21X1 U1437 ( .IN1(n1434), .IN2(n1435), .S(n1436), .Q(n1433) );
  XOR3X1 U1438 ( .IN1(keyinput30), .IN2(N351), .IN3(n1437), .Q(n1436) );
  NOR2X0 U1439 ( .IN1(keyinput14), .IN2(n1438), .QN(n1437) );
  NOR2X0 U1440 ( .IN1(keyinput31), .IN2(n1435), .QN(n1434) );
  XNOR2X1 U1441 ( .IN1(N361), .IN2(N369), .Q(n1435) );
  XNOR3X1 U1442 ( .IN1(n1094), .IN2(N316), .IN3(N308), .Q(n1432) );
  XNOR2X1 U1443 ( .IN1(n1072), .IN2(N293), .Q(n1431) );
  AND3X1 U1444 ( .IN1(n1272), .IN2(n1375), .IN3(n1276), .Q(N6648) );
  AND4X1 U1445 ( .IN1(n1334), .IN2(n931), .IN3(n1378), .IN4(n940), .Q(n1276)
         );
  NOR3X0 U1446 ( .IN1(n1374), .IN2(n1039), .IN3(n1030), .QN(N6646) );
  NAND3X0 U1447 ( .IN1(n1017), .IN2(n1013), .IN3(n1360), .QN(n1030) );
  NAND2X0 U1448 ( .IN1(n1439), .IN2(n1440), .QN(n1013) );
  XNOR2X1 U1449 ( .IN1(keyinput58), .IN2(n1441), .Q(n1439) );
  NAND2X0 U1450 ( .IN1(n1053), .IN2(n1032), .QN(n1374) );
  XNOR2X1 U1451 ( .IN1(n1313), .IN2(keyinput51), .Q(n1032) );
  NOR2X0 U1452 ( .IN1(n1041), .IN2(n1040), .QN(n1053) );
  INVX0 U1453 ( .INP(n1054), .ZN(n1040) );
  XOR2X1 U1454 ( .IN1(n1251), .IN2(keyinput70), .Q(n1054) );
  INVX0 U1455 ( .INP(n1046), .ZN(n1041) );
  NOR4X0 U1456 ( .IN1(n1442), .IN2(n1235), .IN3(n1010), .IN4(n1313), .QN(N6643) );
  MUX21X1 U1457 ( .IN1(N307), .IN2(N302), .S(n1443), .Q(n1313) );
  INVX0 U1458 ( .INP(n1360), .ZN(n1010) );
  NOR2X0 U1459 ( .IN1(n1020), .IN2(n996), .QN(n1360) );
  INVX0 U1460 ( .INP(n1353), .ZN(n1020) );
  NOR2X0 U1461 ( .IN1(n1007), .IN2(n1021), .QN(n1353) );
  NAND2X0 U1462 ( .IN1(n1046), .IN2(n1251), .QN(n1235) );
  INVX0 U1463 ( .INP(n1248), .ZN(n1251) );
  AO21X1 U1464 ( .IN1(n1444), .IN2(n1445), .IN3(n1055), .Q(n1248) );
  NOR2X0 U1465 ( .IN1(n1445), .IN2(n1444), .QN(n1055) );
  INVX0 U1466 ( .INP(n1314), .ZN(n1444) );
  MUX21X1 U1467 ( .IN1(N315), .IN2(N308), .S(n1443), .Q(n1314) );
  NOR2X0 U1468 ( .IN1(n1043), .IN2(n1052), .QN(n1046) );
  NOR2X0 U1469 ( .IN1(n1316), .IN2(N490), .QN(n1052) );
  AND2X1 U1470 ( .IN1(N490), .IN2(n1316), .Q(n1043) );
  MUX21X1 U1471 ( .IN1(N323), .IN2(N316), .S(n1443), .Q(n1316) );
  NAND3X0 U1472 ( .IN1(n1044), .IN2(n1348), .IN3(n1017), .QN(n1442) );
  INVX0 U1473 ( .INP(n1370), .ZN(n1017) );
  INVX0 U1474 ( .INP(n1039), .ZN(n1044) );
  MUX21X1 U1475 ( .IN1(N299), .IN2(N293), .S(n1443), .Q(n1039) );
  AND4X1 U1476 ( .IN1(n962), .IN2(n931), .IN3(n1272), .IN4(n990), .Q(N6641) );
  XNOR2X1 U1477 ( .IN1(n1375), .IN2(keyinput68), .Q(n990) );
  INVX0 U1478 ( .INP(n1267), .ZN(n1375) );
  AO21X1 U1479 ( .IN1(n1307), .IN2(n1446), .IN3(n1377), .Q(n1267) );
  NOR2X0 U1480 ( .IN1(n1307), .IN2(n1446), .QN(n1377) );
  XOR2X1 U1481 ( .IN1(keyinput37), .IN2(n1447), .Q(n1307) );
  MUX21X1 U1482 ( .IN1(N206), .IN2(N209), .S(N335), .Q(n1447) );
  NOR2X0 U1483 ( .IN1(n1278), .IN2(n978), .QN(n1272) );
  INVX0 U1484 ( .INP(n981), .ZN(n978) );
  OA21X1 U1485 ( .IN1(n1304), .IN2(N457), .IN3(n975), .Q(n981) );
  NAND2X0 U1486 ( .IN1(N457), .IN2(n1304), .QN(n975) );
  MUX21X1 U1487 ( .IN1(N210), .IN2(N217), .S(N335), .Q(n1304) );
  NAND2X0 U1488 ( .IN1(n1264), .IN2(n966), .QN(n1278) );
  XOR2X1 U1489 ( .IN1(N468), .IN2(n980), .Q(n966) );
  MUX21X1 U1490 ( .IN1(N218), .IN2(N225), .S(N335), .Q(n980) );
  NOR2X0 U1491 ( .IN1(n971), .IN2(n987), .QN(n1264) );
  NOR2X0 U1492 ( .IN1(n1301), .IN2(N422), .QN(n987) );
  AND2X1 U1493 ( .IN1(N422), .IN2(n1301), .Q(n971) );
  MUX21X1 U1494 ( .IN1(N226), .IN2(N233), .S(N335), .Q(n1301) );
  INVX0 U1495 ( .INP(n922), .ZN(n931) );
  NAND2X0 U1496 ( .IN1(n933), .IN2(n918), .QN(n922) );
  NOR2X0 U1497 ( .IN1(n921), .IN2(n912), .QN(n962) );
  XOR2X1 U1498 ( .IN1(n1378), .IN2(keyinput69), .Q(n912) );
  NAND2X0 U1499 ( .IN1(n940), .IN2(n935), .QN(n921) );
  XNOR2X1 U1500 ( .IN1(keyinput110), .IN2(n1448), .Q(N7515) );
  AOI221X1 U1501 ( .IN1(n851), .IN2(N43), .IN3(n1195), .IN4(n848), .IN5(n1449), 
        .QN(n1448) );
  AO22X1 U1502 ( .IN1(n850), .IN2(N37), .IN3(n1201), .IN4(n847), .Q(n1449) );
  NOR2X0 U1503 ( .IN1(N607), .IN2(N610), .QN(n847) );
  AO222X1 U1504 ( .IN1(N52), .IN2(n1157), .IN3(n1450), .IN4(n855), .IN5(n852), 
        .IN6(n1253), .Q(n1201) );
  XOR2X1 U1505 ( .IN1(n1370), .IN2(n1451), .Q(n1253) );
  OA21X1 U1506 ( .IN1(n1452), .IN2(n1387), .IN3(n1373), .Q(n1451) );
  OR2X1 U1507 ( .IN1(n1090), .IN2(n1326), .Q(n1373) );
  INVX0 U1508 ( .INP(n1348), .ZN(n1387) );
  NAND2X0 U1509 ( .IN1(n1453), .IN2(n1440), .QN(n1348) );
  OR2X1 U1510 ( .IN1(N514), .IN2(n1326), .Q(n1440) );
  XOR2X1 U1511 ( .IN1(n1441), .IN2(keyinput57), .Q(n1453) );
  NAND2X0 U1512 ( .IN1(N514), .IN2(n1326), .QN(n1441) );
  OA21X1 U1513 ( .IN1(n1443), .IN2(N1144), .IN3(n1454), .Q(n1326) );
  OA21X1 U1514 ( .IN1(n1342), .IN2(n1021), .IN3(n1351), .Q(n1452) );
  NAND2X0 U1515 ( .IN1(N523), .IN2(n1325), .QN(n1351) );
  INVX0 U1516 ( .INP(n1019), .ZN(n1021) );
  XOR2X1 U1517 ( .IN1(N523), .IN2(n1325), .Q(n1019) );
  XNOR2X1 U1518 ( .IN1(keyinput39), .IN2(n1455), .Q(n1325) );
  OA22X1 U1519 ( .IN1(n1454), .IN2(n1438), .IN3(N1138), .IN4(n1443), .Q(n1455)
         );
  OA21X1 U1520 ( .IN1(n1007), .IN2(n1366), .IN3(n1023), .Q(n1342) );
  NOR2X0 U1521 ( .IN1(n996), .IN2(N54), .QN(n1366) );
  AO21X1 U1522 ( .IN1(N332), .IN2(N366), .IN3(n1456), .Q(n996) );
  XOR2X1 U1523 ( .IN1(keyinput26), .IN2(n1457), .Q(n1456) );
  NOR2X0 U1524 ( .IN1(n1454), .IN2(n1458), .QN(n1457) );
  INVX0 U1525 ( .INP(N361), .ZN(n1458) );
  INVX0 U1526 ( .INP(n1320), .ZN(n1454) );
  INVX0 U1527 ( .INP(n1018), .ZN(n1007) );
  OA21X1 U1528 ( .IN1(n1322), .IN2(N534), .IN3(n1023), .Q(n1018) );
  NAND2X0 U1529 ( .IN1(N534), .IN2(n1322), .QN(n1023) );
  AO22X1 U1530 ( .IN1(N358), .IN2(N332), .IN3(N351), .IN4(n1320), .Q(n1322) );
  XOR2X1 U1531 ( .IN1(N332), .IN2(keyinput13), .Q(n1320) );
  XNOR2X1 U1532 ( .IN1(n1327), .IN2(N503), .Q(n1370) );
  XOR2X1 U1533 ( .IN1(n1459), .IN2(keyinput40), .Q(n1327) );
  MUX21X1 U1534 ( .IN1(N331), .IN2(N324), .S(n1443), .Q(n1459) );
  INVX0 U1535 ( .INP(N332), .ZN(n1443) );
  AND2X1 U1536 ( .IN1(N607), .IN2(N610), .Q(n850) );
  NOR2X0 U1537 ( .IN1(n1460), .IN2(N607), .QN(n848) );
  AO221X1 U1538 ( .IN1(n1461), .IN2(n855), .IN3(N122), .IN4(n1157), .IN5(n1462), .Q(n1195) );
  XOR2X1 U1539 ( .IN1(n1463), .IN2(keyinput101), .Q(n1462) );
  NAND2X0 U1540 ( .IN1(n1257), .IN2(n852), .QN(n1463) );
  AND2X1 U1541 ( .IN1(N619), .IN2(n907), .Q(n852) );
  XNOR2X1 U1542 ( .IN1(n1378), .IN2(n1464), .Q(n1257) );
  OA21X1 U1543 ( .IN1(n1336), .IN2(n917), .IN3(n1384), .Q(n1464) );
  INVX0 U1544 ( .INP(n940), .ZN(n917) );
  OA21X1 U1545 ( .IN1(n1293), .IN2(N389), .IN3(n1384), .Q(n940) );
  NAND2X0 U1546 ( .IN1(N389), .IN2(n1293), .QN(n1384) );
  XNOR2X1 U1547 ( .IN1(n1465), .IN2(keyinput36), .Q(n1293) );
  AO22X1 U1548 ( .IN1(N264), .IN2(N335), .IN3(N257), .IN4(n1308), .Q(n1465) );
  AOI21X1 U1549 ( .IN1(n1334), .IN2(n1333), .IN3(n1401), .QN(n1336) );
  NOR2X0 U1550 ( .IN1(n875), .IN2(n1292), .QN(n1401) );
  AO21X1 U1551 ( .IN1(n933), .IN2(n1331), .IN3(n1466), .Q(n1333) );
  INVX0 U1552 ( .INP(n1383), .ZN(n1466) );
  AO21X1 U1553 ( .IN1(N4), .IN2(n918), .IN3(n953), .Q(n1331) );
  INVX0 U1554 ( .INP(n1467), .ZN(n953) );
  OA21X1 U1555 ( .IN1(n932), .IN2(N374), .IN3(n1467), .Q(n918) );
  NAND2X0 U1556 ( .IN1(N374), .IN2(n932), .QN(n1467) );
  AO22X1 U1557 ( .IN1(N288), .IN2(N335), .IN3(N281), .IN4(n1308), .Q(n932) );
  OA21X1 U1558 ( .IN1(n1298), .IN2(N411), .IN3(n1383), .Q(n933) );
  NAND2X0 U1559 ( .IN1(N411), .IN2(n1298), .QN(n1383) );
  XNOR2X1 U1560 ( .IN1(n1468), .IN2(keyinput35), .Q(n1298) );
  AO22X1 U1561 ( .IN1(N280), .IN2(N335), .IN3(N273), .IN4(n1308), .Q(n1468) );
  XOR2X1 U1562 ( .IN1(n935), .IN2(keyinput67), .Q(n1334) );
  XOR2X1 U1563 ( .IN1(n1292), .IN2(n875), .Q(n935) );
  AOI22X1 U1564 ( .IN1(N272), .IN2(N335), .IN3(N265), .IN4(n1308), .QN(n1292)
         );
  XOR2X1 U1565 ( .IN1(N335), .IN2(keyinput10), .Q(n1308) );
  XOR2X1 U1566 ( .IN1(N435), .IN2(n1302), .Q(n1378) );
  MUX21X1 U1567 ( .IN1(N234), .IN2(N241), .S(N335), .Q(n1302) );
  NOR2X0 U1568 ( .IN1(n907), .IN2(N619), .QN(n1157) );
  INVX0 U1569 ( .INP(N625), .ZN(n907) );
  NOR2X0 U1570 ( .IN1(N619), .IN2(N625), .QN(n855) );
  AND2X1 U1571 ( .IN1(N607), .IN2(n1460), .Q(n851) );
  INVX0 U1572 ( .INP(N610), .ZN(n1460) );
  NOR4X0 U1573 ( .IN1(n1469), .IN2(n1470), .IN3(n1155), .IN4(n1335), .QN(N5388) );
  MUX41X1 U1574 ( .IN1(n1471), .IN3(n1472), .IN2(N597), .IN4(N598), .S0(N257), 
        .S1(N389), .Q(n1335) );
  MUX41X1 U1575 ( .IN1(n1471), .IN3(n1472), .IN2(N597), .IN4(N598), .S0(N226), 
        .S1(N422), .Q(n1155) );
  OR3X1 U1576 ( .IN1(n902), .IN2(n1158), .IN3(n1160), .Q(n1470) );
  MUX41X1 U1577 ( .IN1(n1471), .IN3(n1472), .IN2(N597), .IN4(N598), .S0(N210), 
        .S1(N457), .Q(n1160) );
  AOI21X1 U1578 ( .IN1(n1473), .IN2(n1474), .IN3(n1475), .QN(n1158) );
  MUX21X1 U1579 ( .IN1(n1476), .IN2(n1477), .S(N468), .Q(n1475) );
  NOR2X0 U1580 ( .IN1(n1478), .IN2(n1474), .QN(n1477) );
  MUX21X1 U1581 ( .IN1(N598), .IN2(N597), .S(n900), .Q(n1478) );
  INVX0 U1582 ( .INP(n1479), .ZN(n1476) );
  MUX21X1 U1583 ( .IN1(n1472), .IN2(n1471), .S(n900), .Q(n1479) );
  INVX0 U1584 ( .INP(keyinput17), .ZN(n1474) );
  NAND3X0 U1585 ( .IN1(n900), .IN2(n1480), .IN3(N468), .QN(n1473) );
  INVX0 U1586 ( .INP(N597), .ZN(n1480) );
  INVX0 U1587 ( .INP(N218), .ZN(n900) );
  MUX41X1 U1588 ( .IN1(n877), .IN3(N242), .IN2(n878), .IN4(N254), .S0(n1446), 
        .S1(n1427), .Q(n902) );
  INVX0 U1589 ( .INP(N206), .ZN(n1427) );
  INVX0 U1590 ( .INP(N446), .ZN(n1446) );
  OR4X1 U1591 ( .IN1(n1481), .IN2(n1364), .IN3(n1461), .IN4(n1330), .Q(n1469)
         );
  MUX41X1 U1592 ( .IN1(n1471), .IN3(n1472), .IN2(N597), .IN4(N598), .S0(N273), 
        .S1(N411), .Q(n1330) );
  MUX21X1 U1593 ( .IN1(n1482), .IN2(n1483), .S(N435), .Q(n1461) );
  OA22X1 U1594 ( .IN1(N597), .IN2(n1484), .IN3(N598), .IN4(n894), .Q(n1483) );
  XNOR2X1 U1595 ( .IN1(N234), .IN2(keyinput8), .Q(n1484) );
  MUX21X1 U1596 ( .IN1(n1472), .IN2(n1471), .S(n894), .Q(n1482) );
  INVX0 U1597 ( .INP(N234), .ZN(n894) );
  MUX41X1 U1598 ( .IN1(n1471), .IN3(n1472), .IN2(N597), .IN4(N598), .S0(N281), 
        .S1(N374), .Q(n1364) );
  XNOR2X1 U1599 ( .IN1(n1332), .IN2(keyinput52), .Q(n1481) );
  MUX21X1 U1600 ( .IN1(n1485), .IN2(n1486), .S(n875), .Q(n1332) );
  INVX0 U1601 ( .INP(N400), .ZN(n875) );
  AO22X1 U1602 ( .IN1(N265), .IN2(n1472), .IN3(n1487), .IN4(n1471), .Q(n1486)
         );
  XNOR2X1 U1603 ( .IN1(keyinput9), .IN2(n879), .Q(n1487) );
  MUX21X1 U1604 ( .IN1(N598), .IN2(N597), .S(n879), .Q(n1485) );
  INVX0 U1605 ( .INP(N265), .ZN(n879) );
  NOR4X0 U1606 ( .IN1(n1488), .IN2(n1489), .IN3(n1365), .IN4(n1450), .QN(N5240) );
  MUX41X1 U1607 ( .IN1(n1472), .IN3(n1471), .IN2(N598), .IN4(N597), .S0(n1094), 
        .S1(N503), .Q(n1450) );
  INVX0 U1608 ( .INP(N324), .ZN(n1094) );
  MUX41X1 U1609 ( .IN1(N597), .IN3(N598), .IN2(n1471), .IN4(n1472), .S0(N351), 
        .S1(n1101), .Q(n1365) );
  INVX0 U1610 ( .INP(N534), .ZN(n1101) );
  OR3X1 U1611 ( .IN1(n1172), .IN2(n1171), .IN3(n1339), .Q(n1489) );
  MUX41X1 U1612 ( .IN1(N598), .IN3(N597), .IN2(n1472), .IN4(n1471), .S0(n1438), 
        .S1(n1097), .Q(n1339) );
  INVX0 U1613 ( .INP(N523), .ZN(n1097) );
  INVX0 U1614 ( .INP(N341), .ZN(n1438) );
  INVX0 U1615 ( .INP(N596), .ZN(n1471) );
  INVX0 U1616 ( .INP(n1084), .ZN(n1171) );
  NAND2X0 U1617 ( .IN1(n1076), .IN2(n1074), .QN(n1084) );
  NAND2X0 U1618 ( .IN1(n1490), .IN2(n1491), .QN(n1074) );
  INVX0 U1619 ( .INP(N490), .ZN(n1491) );
  MUX21X1 U1620 ( .IN1(n888), .IN2(n887), .S(N316), .Q(n1490) );
  NAND2X0 U1621 ( .IN1(n1492), .IN2(N490), .QN(n1076) );
  MUX21X1 U1622 ( .IN1(N251), .IN2(N248), .S(N316), .Q(n1492) );
  AND3X1 U1623 ( .IN1(n1493), .IN2(n1080), .IN3(n1494), .Q(n1172) );
  XOR2X1 U1624 ( .IN1(n1083), .IN2(keyinput11), .Q(n1494) );
  NAND3X0 U1625 ( .IN1(N308), .IN2(N248), .IN3(N479), .QN(n1083) );
  NAND2X0 U1626 ( .IN1(n1495), .IN2(n1445), .QN(n1080) );
  MUX21X1 U1627 ( .IN1(n888), .IN2(n887), .S(N308), .Q(n1495) );
  INVX0 U1628 ( .INP(N242), .ZN(n887) );
  INVX0 U1629 ( .INP(N254), .ZN(n888) );
  XNOR2X1 U1630 ( .IN1(keyinput19), .IN2(n1082), .Q(n1493) );
  OR3X1 U1631 ( .IN1(n878), .IN2(N308), .IN3(n1445), .Q(n1082) );
  INVX0 U1632 ( .INP(N479), .ZN(n1445) );
  OR4X1 U1633 ( .IN1(n1496), .IN2(n1174), .IN3(n1345), .IN4(n1176), .Q(n1488)
         );
  XOR2X1 U1634 ( .IN1(n1070), .IN2(keyinput24), .Q(n1176) );
  MUX21X1 U1635 ( .IN1(N254), .IN2(N242), .S(N293), .Q(n1070) );
  MUX21X1 U1636 ( .IN1(N598), .IN2(n1472), .S(n1090), .Q(n1345) );
  INVX0 U1637 ( .INP(N514), .ZN(n1090) );
  XOR2X1 U1638 ( .IN1(keyinput0), .IN2(N595), .Q(n1472) );
  XOR2X1 U1639 ( .IN1(keyinput38), .IN2(n1497), .Q(n1174) );
  OA21X1 U1640 ( .IN1(n877), .IN2(n1072), .IN3(n1498), .Q(n1497) );
  XOR2X1 U1641 ( .IN1(n1499), .IN2(keyinput18), .Q(n1498) );
  NAND2X0 U1642 ( .IN1(N251), .IN2(n1072), .QN(n1499) );
  INVX0 U1643 ( .INP(N302), .ZN(n1072) );
  XOR2X1 U1644 ( .IN1(n1086), .IN2(keyinput46), .Q(n1496) );
  MUX21X1 U1645 ( .IN1(n878), .IN2(n877), .S(N361), .Q(n1086) );
  INVX0 U1646 ( .INP(N248), .ZN(n877) );
  INVX0 U1647 ( .INP(N251), .ZN(n878) );
  OA21X1 U1648 ( .IN1(N2623), .IN2(n1500), .IN3(N141), .Q(N4740) );
  MUX21X1 U1649 ( .IN1(N80), .IN2(N82), .S(n1501), .Q(n1500) );
  XOR2X1 U1650 ( .IN1(keyinput53), .IN2(n1502), .Q(N4739) );
  OA21X1 U1651 ( .IN1(N2623), .IN2(n1503), .IN3(N141), .Q(n1502) );
  MUX21X1 U1652 ( .IN1(N23), .IN2(N79), .S(n1501), .Q(n1503) );
  OA21X1 U1653 ( .IN1(n1504), .IN2(n1505), .IN3(N141), .Q(N4738) );
  AO21X1 U1654 ( .IN1(N81), .IN2(N588), .IN3(N2623), .Q(n1505) );
  XNOR2X1 U1655 ( .IN1(n1506), .IN2(keyinput43), .Q(n1504) );
  NAND2X0 U1656 ( .IN1(N26), .IN2(n1501), .QN(n1506) );
  OA21X1 U1657 ( .IN1(N2623), .IN2(n1507), .IN3(N141), .Q(N4737) );
  MUX21X1 U1658 ( .IN1(N25), .IN2(N24), .S(n1501), .Q(n1507) );
  XOR2X1 U1659 ( .IN1(n1508), .IN2(keyinput48), .Q(N4279) );
  NAND2X0 U1660 ( .IN1(N83), .IN2(n1509), .QN(n1508) );
  NAND2X0 U1661 ( .IN1(n1510), .IN2(n1509), .QN(N4278) );
  XNOR2X1 U1662 ( .IN1(n1511), .IN2(keyinput34), .Q(n1510) );
  NAND2X0 U1663 ( .IN1(n1511), .IN2(n1509), .QN(N4275) );
  MUX21X1 U1664 ( .IN1(N34), .IN2(N88), .S(n1501), .Q(n1511) );
  XOR2X1 U1665 ( .IN1(n1512), .IN2(keyinput47), .Q(N4272) );
  NAND2X0 U1666 ( .IN1(n1513), .IN2(n1509), .QN(n1512) );
  MUX21X1 U1667 ( .IN1(N87), .IN2(N86), .S(n1501), .Q(n1513) );
  INVX0 U1668 ( .INP(N588), .ZN(n1501) );
  INVX0 U1669 ( .INP(N299), .ZN(N3613) );
  AND2X1 U1670 ( .IN1(N373), .IN2(N1), .Q(N1972) );
  NAND2X0 U1671 ( .IN1(N140), .IN2(n1509), .QN(N2590) );
  INVX0 U1672 ( .INP(N2623), .ZN(n1509) );
  NAND2X0 U1673 ( .IN1(N31), .IN2(N27), .QN(N2623) );
  XOR2X1 U1674 ( .IN1(n1514), .IN2(keyinput3), .Q(N2061) );
  NAND2X0 U1675 ( .IN1(N556), .IN2(N386), .QN(n1514) );
  NAND2X0 U1676 ( .IN1(n1515), .IN2(N27), .QN(N2060) );
  INVX0 U1677 ( .INP(N591), .ZN(n1515) );
  NOR2X0 U1678 ( .IN1(N592), .IN2(n1516), .QN(N2054) );
  INVX0 U1679 ( .INP(N136), .ZN(n1516) );
  XNOR2X1 U1680 ( .IN1(N358), .IN2(keyinput1), .Q(N1145) );
  INVX0 U1681 ( .INP(N559), .ZN(N1155) );
  XNOR2X1 U1682 ( .IN1(keyinput2), .IN2(n1169), .Q(N1154) );
  INVX0 U1683 ( .INP(N245), .ZN(N1152) );
  AND2X1 U1684 ( .IN1(N145), .IN2(N141), .Q(N1147) );
  INVX0 U1685 ( .INP(N338), .ZN(N1144) );
  INVX0 U1686 ( .INP(N549), .ZN(N1141) );
  NOR2X0 U1687 ( .IN1(N1153), .IN2(n1169), .QN(N1140) );
  INVX0 U1688 ( .INP(N562), .ZN(n1169) );
  INVX0 U1689 ( .INP(N552), .ZN(N1153) );
  INVX0 U1690 ( .INP(N366), .ZN(N1139) );
  INVX0 U1691 ( .INP(N348), .ZN(N1138) );
  INVX0 U1692 ( .INP(N545), .ZN(N1137) );
endmodule

