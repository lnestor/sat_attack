
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473;

  XNOR2X1 U292 ( .IN1(keyinput30), .IN2(n262), .Q(G1347) );
  NOR2X0 U293 ( .IN1(n263), .IN2(n264), .QN(n262) );
  XOR2X1 U294 ( .IN1(n265), .IN2(keyinput21), .Q(n264) );
  NAND3X0 U295 ( .IN1(n266), .IN2(G24), .IN3(n267), .QN(n265) );
  OA21X1 U296 ( .IN1(n268), .IN2(n269), .IN3(n270), .Q(n263) );
  XOR2X1 U297 ( .IN1(n271), .IN2(keyinput29), .Q(G1330) );
  MUX21X1 U298 ( .IN1(n272), .IN2(n273), .S(G7), .Q(n271) );
  NOR2X0 U299 ( .IN1(n274), .IN2(n275), .QN(n273) );
  OR2X1 U300 ( .IN1(n275), .IN2(n274), .Q(n272) );
  XNOR2X1 U301 ( .IN1(G32), .IN2(n276), .Q(G1355) );
  NOR2X0 U302 ( .IN1(n268), .IN2(n277), .QN(n276) );
  OA22X1 U303 ( .IN1(n278), .IN2(n279), .IN3(n280), .IN4(n279), .Q(G1352) );
  XNOR2X1 U304 ( .IN1(n281), .IN2(keyinput22), .Q(n279) );
  OR2X1 U305 ( .IN1(n278), .IN2(n280), .Q(n281) );
  NAND2X0 U306 ( .IN1(n282), .IN2(n283), .QN(n278) );
  NOR2X0 U307 ( .IN1(n284), .IN2(n285), .QN(G1351) );
  XOR2X1 U308 ( .IN1(n286), .IN2(keyinput25), .Q(n285) );
  OR3X1 U309 ( .IN1(n268), .IN2(G28), .IN3(n287), .Q(n286) );
  OA21X1 U310 ( .IN1(n268), .IN2(n287), .IN3(G28), .Q(n284) );
  XNOR2X1 U311 ( .IN1(n288), .IN2(n289), .Q(G1349) );
  NAND2X0 U312 ( .IN1(n290), .IN2(n291), .QN(n288) );
  OA21X1 U313 ( .IN1(n292), .IN2(n293), .IN3(n294), .Q(G1348) );
  XOR2X1 U314 ( .IN1(n295), .IN2(keyinput24), .Q(n294) );
  NAND3X0 U315 ( .IN1(n283), .IN2(n293), .IN3(n290), .QN(n295) );
  INVX0 U316 ( .INP(G25), .ZN(n293) );
  NOR2X0 U317 ( .IN1(n296), .IN2(n287), .QN(n292) );
  XOR2X1 U318 ( .IN1(n297), .IN2(G23), .Q(G1346) );
  NAND2X0 U319 ( .IN1(n267), .IN2(n298), .QN(n297) );
  XOR2X1 U320 ( .IN1(n299), .IN2(G22), .Q(G1345) );
  NAND2X0 U321 ( .IN1(n267), .IN2(n291), .QN(n299) );
  XOR2X1 U322 ( .IN1(n300), .IN2(G21), .Q(G1344) );
  NAND2X0 U323 ( .IN1(n267), .IN2(n283), .QN(n300) );
  INVX0 U324 ( .INP(n269), .ZN(n267) );
  NAND3X0 U325 ( .IN1(n301), .IN2(n302), .IN3(n303), .QN(n269) );
  OA21X1 U326 ( .IN1(G20), .IN2(n304), .IN3(n305), .Q(G1343) );
  XOR2X1 U327 ( .IN1(keyinput23), .IN2(n306), .Q(n305) );
  AND2X1 U328 ( .IN1(n304), .IN2(G20), .Q(n306) );
  NAND2X0 U329 ( .IN1(n307), .IN2(n266), .QN(n304) );
  XOR2X1 U330 ( .IN1(n308), .IN2(G19), .Q(G1342) );
  NAND2X0 U331 ( .IN1(n307), .IN2(n298), .QN(n308) );
  XOR2X1 U332 ( .IN1(n309), .IN2(G18), .Q(G1341) );
  NAND2X0 U333 ( .IN1(n307), .IN2(n291), .QN(n309) );
  XOR2X1 U334 ( .IN1(n310), .IN2(G17), .Q(G1340) );
  NAND2X0 U335 ( .IN1(n307), .IN2(n283), .QN(n310) );
  AND3X1 U336 ( .IN1(n301), .IN2(n302), .IN3(n311), .Q(n307) );
  XNOR2X1 U337 ( .IN1(G16), .IN2(n312), .Q(G1339) );
  NOR2X0 U338 ( .IN1(n313), .IN2(n314), .QN(n312) );
  XNOR2X1 U339 ( .IN1(G15), .IN2(n315), .Q(G1338) );
  NOR2X0 U340 ( .IN1(n274), .IN2(n314), .QN(n315) );
  XNOR2X1 U341 ( .IN1(G14), .IN2(n316), .Q(G1337) );
  NOR2X0 U342 ( .IN1(n302), .IN2(n314), .QN(n316) );
  XNOR2X1 U343 ( .IN1(G13), .IN2(n317), .Q(G1336) );
  NOR2X0 U344 ( .IN1(n318), .IN2(n314), .QN(n317) );
  NAND3X0 U345 ( .IN1(n291), .IN2(n296), .IN3(n319), .QN(n314) );
  XOR2X1 U346 ( .IN1(n320), .IN2(G12), .Q(G1335) );
  NAND2X0 U347 ( .IN1(n321), .IN2(n322), .QN(n320) );
  XOR2X1 U348 ( .IN1(n323), .IN2(G11), .Q(G1334) );
  NAND2X0 U349 ( .IN1(n321), .IN2(n324), .QN(n323) );
  XOR2X1 U350 ( .IN1(n325), .IN2(G10), .Q(G1333) );
  NAND2X0 U351 ( .IN1(n321), .IN2(n326), .QN(n325) );
  XOR2X1 U352 ( .IN1(n327), .IN2(G9), .Q(G1332) );
  NAND2X0 U353 ( .IN1(n321), .IN2(n301), .QN(n327) );
  AND4X1 U354 ( .IN1(n268), .IN2(n291), .IN3(n328), .IN4(n329), .Q(n321) );
  NOR2X0 U355 ( .IN1(n330), .IN2(n331), .QN(n329) );
  XNOR2X1 U356 ( .IN1(keyinput18), .IN2(n283), .Q(n331) );
  XNOR2X1 U357 ( .IN1(G8), .IN2(n332), .Q(G1331) );
  NOR2X0 U358 ( .IN1(n313), .IN2(n275), .QN(n332) );
  XNOR2X1 U359 ( .IN1(G6), .IN2(n333), .Q(G1329) );
  NOR2X0 U360 ( .IN1(n275), .IN2(n302), .QN(n333) );
  XNOR2X1 U361 ( .IN1(G5), .IN2(n334), .Q(G1328) );
  NOR2X0 U362 ( .IN1(n318), .IN2(n275), .QN(n334) );
  NAND3X0 U363 ( .IN1(n283), .IN2(n335), .IN3(n319), .QN(n275) );
  AND3X1 U364 ( .IN1(n328), .IN2(n330), .IN3(n266), .Q(n319) );
  XNOR2X1 U365 ( .IN1(G4), .IN2(n336), .Q(G1327) );
  NOR2X0 U366 ( .IN1(n337), .IN2(n313), .QN(n336) );
  MUX21X1 U367 ( .IN1(n338), .IN2(n339), .S(n340), .Q(G1326) );
  NAND2X0 U368 ( .IN1(n341), .IN2(n324), .QN(n339) );
  NOR2X0 U369 ( .IN1(n274), .IN2(n337), .QN(n338) );
  XNOR2X1 U370 ( .IN1(G2), .IN2(n342), .Q(G1325) );
  NOR2X0 U371 ( .IN1(n337), .IN2(n302), .QN(n342) );
  MUX21X1 U372 ( .IN1(n343), .IN2(n344), .S(G1), .Q(G1324) );
  NOR2X0 U373 ( .IN1(n318), .IN2(n337), .QN(n344) );
  INVX0 U374 ( .INP(n341), .ZN(n337) );
  NAND2X0 U375 ( .IN1(n301), .IN2(n341), .QN(n343) );
  XNOR2X1 U376 ( .IN1(n345), .IN2(keyinput20), .Q(n341) );
  NAND4X0 U377 ( .IN1(n335), .IN2(n346), .IN3(n328), .IN4(n268), .QN(n345) );
  INVX0 U378 ( .INP(n266), .ZN(n268) );
  INVX0 U379 ( .INP(n347), .ZN(n328) );
  MUX21X1 U380 ( .IN1(n348), .IN2(n349), .S(n301), .Q(n347) );
  NAND3X0 U381 ( .IN1(n274), .IN2(n302), .IN3(n350), .QN(n349) );
  XNOR2X1 U382 ( .IN1(n313), .IN2(keyinput17), .Q(n350) );
  OA22X1 U383 ( .IN1(n326), .IN2(n351), .IN3(n322), .IN4(n324), .Q(n348) );
  XNOR2X1 U384 ( .IN1(n324), .IN2(n352), .Q(n351) );
  NOR2X0 U385 ( .IN1(keyinput16), .IN2(n313), .QN(n352) );
  INVX0 U386 ( .INP(n318), .ZN(n301) );
  XOR2X1 U387 ( .IN1(n353), .IN2(keyinput28), .Q(G1354) );
  MUX21X1 U388 ( .IN1(n354), .IN2(n355), .S(n356), .Q(n353) );
  NAND2X0 U389 ( .IN1(n282), .IN2(n298), .QN(n355) );
  NOR2X0 U390 ( .IN1(n330), .IN2(n277), .QN(n354) );
  XOR3X1 U391 ( .IN1(keyinput31), .IN2(keyinput27), .IN3(n357), .Q(G1353) );
  MUX21X1 U392 ( .IN1(n358), .IN2(n359), .S(n360), .Q(n357) );
  NAND2X0 U393 ( .IN1(n282), .IN2(n291), .QN(n359) );
  INVX0 U394 ( .INP(n277), .ZN(n282) );
  NOR2X0 U395 ( .IN1(n335), .IN2(n277), .QN(n358) );
  NAND3X0 U396 ( .IN1(n303), .IN2(n318), .IN3(n326), .QN(n277) );
  AND3X1 U397 ( .IN1(n322), .IN2(n361), .IN3(n274), .Q(n303) );
  INVX0 U398 ( .INP(n324), .ZN(n274) );
  XOR2X1 U399 ( .IN1(n362), .IN2(keyinput26), .Q(G1350) );
  MUX21X1 U400 ( .IN1(n363), .IN2(n364), .S(G27), .Q(n362) );
  NOR2X0 U401 ( .IN1(n330), .IN2(n287), .QN(n364) );
  NAND2X0 U402 ( .IN1(n290), .IN2(n298), .QN(n363) );
  INVX0 U403 ( .INP(n330), .ZN(n298) );
  INVX0 U404 ( .INP(n287), .ZN(n290) );
  NAND3X0 U405 ( .IN1(n326), .IN2(n318), .IN3(n311), .QN(n287) );
  AND3X1 U406 ( .IN1(n324), .IN2(n361), .IN3(n313), .Q(n311) );
  INVX0 U407 ( .INP(n322), .ZN(n313) );
  MUX21X1 U408 ( .IN1(n365), .IN2(n366), .S(n367), .Q(n322) );
  XOR3X1 U409 ( .IN1(G16), .IN2(G12), .IN3(n368), .Q(n367) );
  XNOR3X1 U410 ( .IN1(keyinput5), .IN2(n369), .IN3(G4), .Q(n368) );
  INVX0 U411 ( .INP(G8), .ZN(n369) );
  AND2X1 U412 ( .IN1(n370), .IN2(n371), .Q(n366) );
  NAND2X0 U413 ( .IN1(n371), .IN2(n370), .QN(n365) );
  AO21X1 U414 ( .IN1(G36), .IN2(G41), .IN3(n372), .Q(n370) );
  NAND3X0 U415 ( .IN1(G36), .IN2(G41), .IN3(n372), .QN(n371) );
  XOR2X1 U416 ( .IN1(n373), .IN2(n374), .Q(n372) );
  NAND2X0 U417 ( .IN1(n375), .IN2(n376), .QN(n361) );
  OR3X1 U418 ( .IN1(n266), .IN2(n346), .IN3(n291), .Q(n376) );
  NOR2X0 U419 ( .IN1(n330), .IN2(n296), .QN(n346) );
  NAND3X0 U420 ( .IN1(n377), .IN2(n330), .IN3(n296), .QN(n375) );
  INVX0 U421 ( .INP(n283), .ZN(n296) );
  MUX21X1 U422 ( .IN1(n378), .IN2(n379), .S(n380), .Q(n283) );
  XOR3X1 U423 ( .IN1(G21), .IN2(G17), .IN3(n381), .Q(n380) );
  XNOR2X1 U424 ( .IN1(n280), .IN2(G25), .Q(n381) );
  INVX0 U425 ( .INP(G29), .ZN(n280) );
  NAND2X0 U426 ( .IN1(n382), .IN2(n383), .QN(n379) );
  AND2X1 U427 ( .IN1(n383), .IN2(n382), .Q(n378) );
  NAND3X0 U428 ( .IN1(G37), .IN2(G41), .IN3(n384), .QN(n382) );
  AO21X1 U429 ( .IN1(G37), .IN2(G41), .IN3(n384), .Q(n383) );
  XNOR2X1 U430 ( .IN1(n385), .IN2(n386), .Q(n384) );
  AO22X1 U431 ( .IN1(n387), .IN2(n388), .IN3(n389), .IN4(n390), .Q(n330) );
  XOR2X1 U432 ( .IN1(n391), .IN2(keyinput13), .Q(n390) );
  AND2X1 U433 ( .IN1(n392), .IN2(n393), .Q(n389) );
  NAND2X0 U434 ( .IN1(n393), .IN2(n392), .QN(n388) );
  AO21X1 U435 ( .IN1(G41), .IN2(G39), .IN3(n394), .Q(n392) );
  NAND3X0 U436 ( .IN1(G41), .IN2(G39), .IN3(n394), .QN(n393) );
  XNOR2X1 U437 ( .IN1(n395), .IN2(n386), .Q(n394) );
  XOR3X1 U438 ( .IN1(G2), .IN2(n396), .IN3(G1), .Q(n386) );
  OA21X1 U439 ( .IN1(G4), .IN2(n340), .IN3(n397), .Q(n396) );
  XOR2X1 U440 ( .IN1(n398), .IN2(keyinput2), .Q(n397) );
  NAND2X0 U441 ( .IN1(G4), .IN2(n340), .QN(n398) );
  XNOR2X1 U442 ( .IN1(keyinput13), .IN2(n391), .Q(n387) );
  AO21X1 U443 ( .IN1(n399), .IN2(n400), .IN3(n401), .Q(n391) );
  XOR2X1 U444 ( .IN1(n402), .IN2(keyinput12), .Q(n401) );
  NAND2X0 U445 ( .IN1(n403), .IN2(n400), .QN(n402) );
  NAND2X0 U446 ( .IN1(n399), .IN2(n403), .QN(n400) );
  AO21X1 U447 ( .IN1(G27), .IN2(n356), .IN3(n404), .Q(n403) );
  XOR2X1 U448 ( .IN1(n405), .IN2(keyinput3), .Q(n404) );
  OR2X1 U449 ( .IN1(n356), .IN2(G27), .Q(n405) );
  INVX0 U450 ( .INP(G31), .ZN(n356) );
  XOR2X1 U451 ( .IN1(G23), .IN2(G19), .Q(n399) );
  NAND2X0 U452 ( .IN1(n266), .IN2(n406), .QN(n377) );
  XNOR2X1 U453 ( .IN1(keyinput19), .IN2(n335), .Q(n406) );
  INVX0 U454 ( .INP(n291), .ZN(n335) );
  XOR3X1 U455 ( .IN1(n407), .IN2(n408), .IN3(n409), .Q(n291) );
  XOR3X1 U456 ( .IN1(keyinput0), .IN2(n410), .IN3(n411), .Q(n409) );
  NAND2X0 U457 ( .IN1(G38), .IN2(G41), .QN(n411) );
  OA21X1 U458 ( .IN1(n412), .IN2(n413), .IN3(n414), .Q(n410) );
  XOR2X1 U459 ( .IN1(n415), .IN2(keyinput11), .Q(n414) );
  NAND2X0 U460 ( .IN1(n412), .IN2(n413), .QN(n415) );
  XOR3X1 U461 ( .IN1(keyinput6), .IN2(G22), .IN3(G18), .Q(n413) );
  AOI21X1 U462 ( .IN1(n289), .IN2(n360), .IN3(n416), .QN(n412) );
  XOR2X1 U463 ( .IN1(keyinput1), .IN2(n417), .Q(n416) );
  NOR2X0 U464 ( .IN1(n289), .IN2(n360), .QN(n417) );
  INVX0 U465 ( .INP(G30), .ZN(n360) );
  INVX0 U466 ( .INP(G26), .ZN(n289) );
  INVX0 U467 ( .INP(n395), .ZN(n408) );
  XNOR3X1 U468 ( .IN1(G11), .IN2(G10), .IN3(n418), .Q(n395) );
  XNOR2X1 U469 ( .IN1(G12), .IN2(G9), .Q(n418) );
  MUX21X1 U470 ( .IN1(n419), .IN2(n420), .S(n421), .Q(n266) );
  XNOR3X1 U471 ( .IN1(n270), .IN2(G20), .IN3(n422), .Q(n421) );
  XOR2X1 U472 ( .IN1(G32), .IN2(G28), .Q(n422) );
  INVX0 U473 ( .INP(G24), .ZN(n270) );
  NAND2X0 U474 ( .IN1(n423), .IN2(n424), .QN(n420) );
  AND2X1 U475 ( .IN1(n424), .IN2(n423), .Q(n419) );
  NAND3X0 U476 ( .IN1(G41), .IN2(n425), .IN3(G40), .QN(n423) );
  AO21X1 U477 ( .IN1(G40), .IN2(G41), .IN3(n425), .Q(n424) );
  XOR2X1 U478 ( .IN1(n407), .IN2(n385), .Q(n425) );
  XOR3X1 U479 ( .IN1(n426), .IN2(G5), .IN3(n427), .Q(n385) );
  XNOR2X1 U480 ( .IN1(G7), .IN2(G8), .Q(n427) );
  XNOR3X1 U481 ( .IN1(G14), .IN2(G13), .IN3(n428), .Q(n407) );
  XNOR2X1 U482 ( .IN1(G15), .IN2(G16), .Q(n428) );
  XNOR3X1 U483 ( .IN1(n429), .IN2(n430), .IN3(n431), .Q(n324) );
  MUX21X1 U484 ( .IN1(n432), .IN2(n433), .S(n434), .Q(n431) );
  OA21X1 U485 ( .IN1(n435), .IN2(n436), .IN3(n437), .Q(n434) );
  XOR2X1 U486 ( .IN1(n438), .IN2(keyinput14), .Q(n437) );
  NAND2X0 U487 ( .IN1(n435), .IN2(n436), .QN(n438) );
  AND2X1 U488 ( .IN1(G41), .IN2(G35), .Q(n433) );
  NAND2X0 U489 ( .IN1(G35), .IN2(G41), .QN(n432) );
  XNOR3X1 U490 ( .IN1(keyinput4), .IN2(G7), .IN3(n340), .Q(n430) );
  INVX0 U491 ( .INP(G3), .ZN(n340) );
  XNOR2X1 U492 ( .IN1(n439), .IN2(G11), .Q(n429) );
  INVX0 U493 ( .INP(G15), .ZN(n439) );
  XNOR3X1 U494 ( .IN1(G1), .IN2(n440), .IN3(n441), .Q(n318) );
  NAND2X0 U495 ( .IN1(n442), .IN2(n443), .QN(n441) );
  NAND3X0 U496 ( .IN1(G41), .IN2(n444), .IN3(G33), .QN(n443) );
  XOR2X1 U497 ( .IN1(keyinput15), .IN2(n445), .Q(n442) );
  NOR2X0 U498 ( .IN1(n446), .IN2(n447), .QN(n445) );
  XOR2X1 U499 ( .IN1(n436), .IN2(n373), .Q(n447) );
  INVX0 U500 ( .INP(n444), .ZN(n446) );
  NAND3X0 U501 ( .IN1(G33), .IN2(G41), .IN3(n448), .QN(n444) );
  XNOR2X1 U502 ( .IN1(n436), .IN2(n373), .Q(n448) );
  AO21X1 U503 ( .IN1(n449), .IN2(n450), .IN3(n451), .Q(n373) );
  XOR2X1 U504 ( .IN1(keyinput9), .IN2(n452), .Q(n451) );
  NOR2X0 U505 ( .IN1(n449), .IN2(n450), .QN(n452) );
  XOR2X1 U506 ( .IN1(G23), .IN2(G24), .Q(n450) );
  XNOR2X1 U507 ( .IN1(G21), .IN2(G22), .Q(n449) );
  AO21X1 U508 ( .IN1(n453), .IN2(n454), .IN3(n455), .Q(n436) );
  XOR2X1 U509 ( .IN1(n456), .IN2(keyinput7), .Q(n455) );
  NAND2X0 U510 ( .IN1(n457), .IN2(n458), .QN(n456) );
  XOR2X1 U511 ( .IN1(G18), .IN2(G17), .Q(n458) );
  XOR2X1 U512 ( .IN1(G20), .IN2(G19), .Q(n457) );
  XNOR2X1 U513 ( .IN1(G17), .IN2(G18), .Q(n454) );
  XNOR2X1 U514 ( .IN1(G19), .IN2(G20), .Q(n453) );
  XOR3X1 U515 ( .IN1(G9), .IN2(G5), .IN3(G13), .Q(n440) );
  INVX0 U516 ( .INP(n302), .ZN(n326) );
  XNOR3X1 U517 ( .IN1(n459), .IN2(n435), .IN3(n460), .Q(n302) );
  XOR2X1 U518 ( .IN1(n461), .IN2(n374), .Q(n460) );
  AOI21X1 U519 ( .IN1(n462), .IN2(n463), .IN3(n464), .QN(n374) );
  XOR2X1 U520 ( .IN1(keyinput8), .IN2(n465), .Q(n464) );
  NOR2X0 U521 ( .IN1(n462), .IN2(n463), .QN(n465) );
  XNOR2X1 U522 ( .IN1(G32), .IN2(G31), .Q(n463) );
  XNOR2X1 U523 ( .IN1(G29), .IN2(G30), .Q(n462) );
  NAND2X0 U524 ( .IN1(G34), .IN2(G41), .QN(n461) );
  XNOR3X1 U525 ( .IN1(G26), .IN2(G25), .IN3(n466), .Q(n435) );
  XNOR2X1 U526 ( .IN1(G27), .IN2(G28), .Q(n466) );
  OA21X1 U527 ( .IN1(n467), .IN2(n468), .IN3(n469), .Q(n459) );
  XOR2X1 U528 ( .IN1(keyinput10), .IN2(n470), .Q(n469) );
  NOR2X0 U529 ( .IN1(n471), .IN2(n472), .QN(n470) );
  XNOR2X1 U530 ( .IN1(n426), .IN2(G2), .Q(n472) );
  INVX0 U531 ( .INP(G6), .ZN(n426) );
  XNOR2X1 U532 ( .IN1(G10), .IN2(G14), .Q(n471) );
  XNOR2X1 U533 ( .IN1(n473), .IN2(G10), .Q(n468) );
  INVX0 U534 ( .INP(G14), .ZN(n473) );
  XNOR2X1 U535 ( .IN1(G2), .IN2(G6), .Q(n467) );
endmodule

