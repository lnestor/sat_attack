
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550;

  XOR2X1 U339 ( .IN1(n307), .IN2(G32), .Q(G1355) );
  NAND2X0 U340 ( .IN1(n308), .IN2(n309), .QN(n307) );
  XOR2X1 U341 ( .IN1(n310), .IN2(G31), .Q(G1354) );
  NAND2X0 U342 ( .IN1(n308), .IN2(n311), .QN(n310) );
  XOR2X1 U343 ( .IN1(n312), .IN2(G30), .Q(G1353) );
  NAND2X0 U344 ( .IN1(n308), .IN2(n313), .QN(n312) );
  XOR2X1 U345 ( .IN1(n314), .IN2(G29), .Q(G1352) );
  NAND2X0 U346 ( .IN1(n308), .IN2(n315), .QN(n314) );
  AND4X1 U347 ( .IN1(n316), .IN2(n317), .IN3(n318), .IN4(n319), .Q(n308) );
  XNOR2X1 U348 ( .IN1(G28), .IN2(n320), .Q(G1351) );
  NOR2X0 U349 ( .IN1(n321), .IN2(n322), .QN(n320) );
  XNOR2X1 U350 ( .IN1(G27), .IN2(n323), .Q(G1350) );
  NOR2X0 U351 ( .IN1(n324), .IN2(n322), .QN(n323) );
  XNOR2X1 U352 ( .IN1(G26), .IN2(n325), .Q(G1349) );
  NOR2X0 U353 ( .IN1(n326), .IN2(n322), .QN(n325) );
  XNOR2X1 U354 ( .IN1(G25), .IN2(n327), .Q(G1348) );
  NOR2X0 U355 ( .IN1(n328), .IN2(n322), .QN(n327) );
  NAND4X0 U356 ( .IN1(n329), .IN2(n319), .IN3(n318), .IN4(n330), .QN(n322) );
  NOR2X0 U357 ( .IN1(n331), .IN2(n317), .QN(n330) );
  XNOR2X1 U358 ( .IN1(G24), .IN2(n332), .Q(G1347) );
  NOR2X0 U359 ( .IN1(n321), .IN2(n333), .QN(n332) );
  XNOR2X1 U360 ( .IN1(G23), .IN2(n334), .Q(G1346) );
  NOR2X0 U361 ( .IN1(n324), .IN2(n333), .QN(n334) );
  XNOR2X1 U362 ( .IN1(G22), .IN2(n335), .Q(G1345) );
  NOR2X0 U363 ( .IN1(n326), .IN2(n333), .QN(n335) );
  XNOR2X1 U364 ( .IN1(G21), .IN2(n336), .Q(G1344) );
  NOR2X0 U365 ( .IN1(n328), .IN2(n333), .QN(n336) );
  NAND4X0 U366 ( .IN1(n331), .IN2(n319), .IN3(n317), .IN4(n337), .QN(n333) );
  NOR2X0 U367 ( .IN1(n318), .IN2(n329), .QN(n337) );
  XOR2X1 U368 ( .IN1(n338), .IN2(G20), .Q(G1343) );
  NAND2X0 U369 ( .IN1(n339), .IN2(n309), .QN(n338) );
  XOR2X1 U370 ( .IN1(n340), .IN2(G19), .Q(G1342) );
  NAND2X0 U371 ( .IN1(n339), .IN2(n311), .QN(n340) );
  XOR2X1 U372 ( .IN1(n341), .IN2(G18), .Q(G1341) );
  NAND2X0 U373 ( .IN1(n339), .IN2(n313), .QN(n341) );
  XOR2X1 U374 ( .IN1(n342), .IN2(G17), .Q(G1340) );
  NAND2X0 U375 ( .IN1(n339), .IN2(n315), .QN(n342) );
  AND4X1 U376 ( .IN1(n343), .IN2(n329), .IN3(n331), .IN4(n319), .Q(n339) );
  NAND2X0 U377 ( .IN1(n344), .IN2(n345), .QN(n319) );
  OR3X1 U378 ( .IN1(n313), .IN2(n346), .IN3(n309), .Q(n345) );
  OR3X1 U379 ( .IN1(n311), .IN2(n347), .IN3(n315), .Q(n344) );
  XOR2X1 U380 ( .IN1(n348), .IN2(G16), .Q(G1339) );
  NAND2X0 U381 ( .IN1(n349), .IN2(n350), .QN(n348) );
  XNOR2X1 U382 ( .IN1(n351), .IN2(n352), .Q(G1338) );
  NAND2X0 U383 ( .IN1(n349), .IN2(n353), .QN(n351) );
  XOR2X1 U384 ( .IN1(n354), .IN2(G14), .Q(G1337) );
  NAND2X0 U385 ( .IN1(n349), .IN2(n355), .QN(n354) );
  XOR2X1 U386 ( .IN1(n356), .IN2(G13), .Q(G1336) );
  NAND2X0 U387 ( .IN1(n349), .IN2(n357), .QN(n356) );
  AND4X1 U388 ( .IN1(n347), .IN2(n328), .IN3(n324), .IN4(n358), .Q(n349) );
  NOR2X0 U389 ( .IN1(n326), .IN2(n321), .QN(n347) );
  XNOR2X1 U390 ( .IN1(G12), .IN2(n359), .Q(G1335) );
  NOR2X0 U391 ( .IN1(n329), .IN2(n360), .QN(n359) );
  XNOR2X1 U392 ( .IN1(G11), .IN2(n361), .Q(G1334) );
  NOR2X0 U393 ( .IN1(n317), .IN2(n360), .QN(n361) );
  XNOR2X1 U394 ( .IN1(G10), .IN2(n362), .Q(G1333) );
  NOR2X0 U395 ( .IN1(n331), .IN2(n360), .QN(n362) );
  XNOR2X1 U396 ( .IN1(G9), .IN2(n363), .Q(G1332) );
  NOR2X0 U397 ( .IN1(n318), .IN2(n360), .QN(n363) );
  NAND4X0 U398 ( .IN1(n328), .IN2(n358), .IN3(n321), .IN4(n364), .QN(n360) );
  NOR2X0 U399 ( .IN1(n324), .IN2(n326), .QN(n364) );
  XNOR2X1 U400 ( .IN1(G8), .IN2(n365), .Q(G1331) );
  NOR2X0 U401 ( .IN1(n329), .IN2(n366), .QN(n365) );
  XNOR2X1 U402 ( .IN1(G7), .IN2(n367), .Q(G1330) );
  NOR2X0 U403 ( .IN1(n317), .IN2(n366), .QN(n367) );
  XNOR2X1 U404 ( .IN1(G6), .IN2(n368), .Q(G1329) );
  NOR2X0 U405 ( .IN1(n331), .IN2(n366), .QN(n368) );
  XNOR2X1 U406 ( .IN1(G5), .IN2(n369), .Q(G1328) );
  NOR2X0 U407 ( .IN1(n318), .IN2(n366), .QN(n369) );
  NAND4X0 U408 ( .IN1(n324), .IN2(n358), .IN3(n326), .IN4(n370), .QN(n366) );
  NOR2X0 U409 ( .IN1(n321), .IN2(n328), .QN(n370) );
  XOR2X1 U410 ( .IN1(n371), .IN2(G4), .Q(G1327) );
  NAND2X0 U411 ( .IN1(n372), .IN2(n350), .QN(n371) );
  XOR2X1 U412 ( .IN1(n373), .IN2(G3), .Q(G1326) );
  NAND2X0 U413 ( .IN1(n372), .IN2(n353), .QN(n373) );
  XOR2X1 U414 ( .IN1(n374), .IN2(G2), .Q(G1325) );
  NAND2X0 U415 ( .IN1(n372), .IN2(n355), .QN(n374) );
  XOR2X1 U416 ( .IN1(n375), .IN2(G1), .Q(G1324) );
  NAND2X0 U417 ( .IN1(n372), .IN2(n357), .QN(n375) );
  AND4X1 U418 ( .IN1(n346), .IN2(n321), .IN3(n326), .IN4(n358), .Q(n372) );
  NAND2X0 U419 ( .IN1(n376), .IN2(n377), .QN(n358) );
  OR3X1 U420 ( .IN1(n355), .IN2(n343), .IN3(n350), .Q(n377) );
  NOR2X0 U421 ( .IN1(n318), .IN2(n317), .QN(n343) );
  INVX0 U422 ( .INP(n353), .ZN(n317) );
  INVX0 U423 ( .INP(n357), .ZN(n318) );
  INVX0 U424 ( .INP(n331), .ZN(n355) );
  OR3X1 U425 ( .IN1(n357), .IN2(n316), .IN3(n353), .Q(n376) );
  MUX21X1 U426 ( .IN1(n378), .IN2(n379), .S(n380), .Q(n353) );
  XNOR3X1 U427 ( .IN1(n352), .IN2(G11), .IN3(n381), .Q(n380) );
  XOR2X1 U428 ( .IN1(G7), .IN2(G3), .Q(n381) );
  INVX0 U429 ( .INP(G15), .ZN(n352) );
  XOR2X1 U430 ( .IN1(n382), .IN2(n383), .Q(n379) );
  XNOR2X1 U431 ( .IN1(n382), .IN2(n383), .Q(n378) );
  AND2X1 U432 ( .IN1(G35), .IN2(G41), .Q(n383) );
  OA21X1 U433 ( .IN1(n384), .IN2(n385), .IN3(n386), .Q(n382) );
  XNOR2X1 U434 ( .IN1(keyinput61), .IN2(n387), .Q(n386) );
  NOR2X0 U435 ( .IN1(n388), .IN2(n384), .QN(n387) );
  XNOR2X1 U436 ( .IN1(n389), .IN2(keyinput54), .Q(n384) );
  NAND2X0 U437 ( .IN1(n390), .IN2(n391), .QN(n389) );
  NOR2X0 U438 ( .IN1(n331), .IN2(n329), .QN(n316) );
  INVX0 U439 ( .INP(n350), .ZN(n329) );
  MUX21X1 U440 ( .IN1(n392), .IN2(n393), .S(n394), .Q(n350) );
  XOR3X1 U441 ( .IN1(G16), .IN2(G12), .IN3(n395), .Q(n394) );
  XOR2X1 U442 ( .IN1(G8), .IN2(G4), .Q(n395) );
  XNOR2X1 U443 ( .IN1(n396), .IN2(n397), .Q(n393) );
  XOR2X1 U444 ( .IN1(n397), .IN2(n396), .Q(n392) );
  AND2X1 U445 ( .IN1(n398), .IN2(n399), .Q(n396) );
  XOR2X1 U446 ( .IN1(keyinput62), .IN2(n400), .Q(n399) );
  NOR2X0 U447 ( .IN1(n401), .IN2(n402), .QN(n400) );
  XOR2X1 U448 ( .IN1(keyinput63), .IN2(n403), .Q(n398) );
  NOR2X0 U449 ( .IN1(n404), .IN2(n402), .QN(n403) );
  XNOR2X1 U450 ( .IN1(n405), .IN2(keyinput55), .Q(n402) );
  NAND2X0 U451 ( .IN1(n406), .IN2(n407), .QN(n405) );
  NAND2X0 U452 ( .IN1(G36), .IN2(G41), .QN(n397) );
  XNOR3X1 U453 ( .IN1(G10), .IN2(n408), .IN3(n409), .Q(n331) );
  MUX21X1 U454 ( .IN1(n410), .IN2(n411), .S(n412), .Q(n409) );
  OA21X1 U455 ( .IN1(n385), .IN2(n413), .IN3(n414), .Q(n412) );
  XOR2X1 U456 ( .IN1(n415), .IN2(keyinput60), .Q(n414) );
  OR2X1 U457 ( .IN1(n413), .IN2(n404), .Q(n415) );
  XNOR2X1 U458 ( .IN1(n416), .IN2(keyinput53), .Q(n413) );
  NAND2X0 U459 ( .IN1(n391), .IN2(n407), .QN(n416) );
  INVX0 U460 ( .INP(n404), .ZN(n407) );
  XNOR2X1 U461 ( .IN1(n417), .IN2(keyinput47), .Q(n404) );
  NAND2X0 U462 ( .IN1(n418), .IN2(n419), .QN(n417) );
  XOR2X1 U463 ( .IN1(keyinput39), .IN2(n420), .Q(n419) );
  AND2X1 U464 ( .IN1(n421), .IN2(n422), .Q(n420) );
  XOR2X1 U465 ( .IN1(n423), .IN2(keyinput38), .Q(n418) );
  NAND2X0 U466 ( .IN1(n422), .IN2(n424), .QN(n423) );
  XOR2X1 U467 ( .IN1(n425), .IN2(keyinput23), .Q(n422) );
  NAND2X0 U468 ( .IN1(n424), .IN2(n421), .QN(n425) );
  XNOR3X1 U469 ( .IN1(keyinput15), .IN2(G32), .IN3(G31), .Q(n421) );
  XNOR3X1 U470 ( .IN1(keyinput14), .IN2(G30), .IN3(G29), .Q(n424) );
  INVX0 U471 ( .INP(n385), .ZN(n391) );
  XNOR2X1 U472 ( .IN1(n426), .IN2(keyinput46), .Q(n385) );
  NAND2X0 U473 ( .IN1(n427), .IN2(n428), .QN(n426) );
  XOR2X1 U474 ( .IN1(n429), .IN2(keyinput36), .Q(n428) );
  NAND2X0 U475 ( .IN1(n430), .IN2(n431), .QN(n429) );
  XOR2X1 U476 ( .IN1(n432), .IN2(keyinput37), .Q(n427) );
  NAND2X0 U477 ( .IN1(n433), .IN2(n431), .QN(n432) );
  XNOR2X1 U478 ( .IN1(n434), .IN2(keyinput22), .Q(n431) );
  NAND2X0 U479 ( .IN1(n430), .IN2(n433), .QN(n434) );
  XNOR3X1 U480 ( .IN1(keyinput12), .IN2(G26), .IN3(G25), .Q(n430) );
  XNOR3X1 U481 ( .IN1(keyinput13), .IN2(G28), .IN3(G27), .Q(n433) );
  AND2X1 U482 ( .IN1(G41), .IN2(G34), .Q(n411) );
  NAND2X0 U483 ( .IN1(G34), .IN2(G41), .QN(n410) );
  XOR3X1 U484 ( .IN1(G6), .IN2(G2), .IN3(G14), .Q(n408) );
  MUX21X1 U485 ( .IN1(n435), .IN2(n436), .S(n437), .Q(n357) );
  XOR3X1 U486 ( .IN1(G13), .IN2(G1), .IN3(n438), .Q(n437) );
  XOR2X1 U487 ( .IN1(G9), .IN2(G5), .Q(n438) );
  NAND2X0 U488 ( .IN1(n439), .IN2(n440), .QN(n436) );
  AND2X1 U489 ( .IN1(n440), .IN2(n439), .Q(n435) );
  NAND4X0 U490 ( .IN1(n441), .IN2(G33), .IN3(G41), .IN4(n442), .QN(n439) );
  AO22X1 U491 ( .IN1(G33), .IN2(G41), .IN3(n441), .IN4(n442), .Q(n440) );
  NAND2X0 U492 ( .IN1(n388), .IN2(n401), .QN(n442) );
  XOR2X1 U493 ( .IN1(n443), .IN2(keyinput52), .Q(n441) );
  NAND2X0 U494 ( .IN1(n390), .IN2(n406), .QN(n443) );
  INVX0 U495 ( .INP(n401), .ZN(n406) );
  XNOR2X1 U496 ( .IN1(n444), .IN2(keyinput45), .Q(n401) );
  NAND2X0 U497 ( .IN1(n445), .IN2(n446), .QN(n444) );
  XOR2X1 U498 ( .IN1(keyinput34), .IN2(n447), .Q(n446) );
  NOR2X0 U499 ( .IN1(n448), .IN2(n449), .QN(n447) );
  XOR2X1 U500 ( .IN1(keyinput35), .IN2(n450), .Q(n445) );
  NOR2X0 U501 ( .IN1(n451), .IN2(n449), .QN(n450) );
  XNOR2X1 U502 ( .IN1(n452), .IN2(keyinput21), .Q(n449) );
  OR2X1 U503 ( .IN1(n448), .IN2(n451), .Q(n452) );
  XOR3X1 U504 ( .IN1(keyinput10), .IN2(G22), .IN3(G21), .Q(n448) );
  XNOR3X1 U505 ( .IN1(keyinput11), .IN2(G24), .IN3(G23), .Q(n451) );
  INVX0 U506 ( .INP(n388), .ZN(n390) );
  XNOR2X1 U507 ( .IN1(n453), .IN2(keyinput44), .Q(n388) );
  NAND2X0 U508 ( .IN1(n454), .IN2(n455), .QN(n453) );
  XOR2X1 U509 ( .IN1(n456), .IN2(keyinput32), .Q(n455) );
  NAND2X0 U510 ( .IN1(n457), .IN2(n458), .QN(n456) );
  XOR2X1 U511 ( .IN1(n459), .IN2(keyinput33), .Q(n454) );
  NAND2X0 U512 ( .IN1(n460), .IN2(n458), .QN(n459) );
  XNOR2X1 U513 ( .IN1(n461), .IN2(keyinput20), .Q(n458) );
  NAND2X0 U514 ( .IN1(n457), .IN2(n460), .QN(n461) );
  XNOR3X1 U515 ( .IN1(keyinput8), .IN2(G18), .IN3(G17), .Q(n457) );
  XNOR3X1 U516 ( .IN1(keyinput9), .IN2(G20), .IN3(G19), .Q(n460) );
  INVX0 U517 ( .INP(n313), .ZN(n326) );
  MUX21X1 U518 ( .IN1(n462), .IN2(n463), .S(n464), .Q(n313) );
  XOR3X1 U519 ( .IN1(G22), .IN2(G18), .IN3(n465), .Q(n464) );
  XOR2X1 U520 ( .IN1(G30), .IN2(G26), .Q(n465) );
  XNOR2X1 U521 ( .IN1(n466), .IN2(n467), .Q(n463) );
  XOR2X1 U522 ( .IN1(n466), .IN2(n467), .Q(n462) );
  AND2X1 U523 ( .IN1(G38), .IN2(G41), .Q(n467) );
  NAND2X0 U524 ( .IN1(n468), .IN2(n469), .QN(n466) );
  XOR2X1 U525 ( .IN1(keyinput59), .IN2(n470), .Q(n469) );
  NOR2X0 U526 ( .IN1(n471), .IN2(n472), .QN(n470) );
  XOR2X1 U527 ( .IN1(n473), .IN2(keyinput58), .Q(n468) );
  OR2X1 U528 ( .IN1(n472), .IN2(n474), .Q(n473) );
  XNOR2X1 U529 ( .IN1(n475), .IN2(keyinput49), .Q(n472) );
  NAND2X0 U530 ( .IN1(n476), .IN2(n477), .QN(n475) );
  INVX0 U531 ( .INP(n309), .ZN(n321) );
  MUX21X1 U532 ( .IN1(n478), .IN2(n479), .S(n480), .Q(n309) );
  XNOR3X1 U533 ( .IN1(n481), .IN2(G20), .IN3(n482), .Q(n480) );
  XOR2X1 U534 ( .IN1(G32), .IN2(G28), .Q(n482) );
  INVX0 U535 ( .INP(G24), .ZN(n481) );
  NAND2X0 U536 ( .IN1(n483), .IN2(n484), .QN(n479) );
  AND2X1 U537 ( .IN1(n484), .IN2(n483), .Q(n478) );
  NAND4X0 U538 ( .IN1(n485), .IN2(G40), .IN3(G41), .IN4(n486), .QN(n483) );
  AO22X1 U539 ( .IN1(G40), .IN2(G41), .IN3(n485), .IN4(n486), .Q(n484) );
  NAND2X0 U540 ( .IN1(n471), .IN2(n487), .QN(n486) );
  INVX0 U541 ( .INP(n476), .ZN(n471) );
  XOR2X1 U542 ( .IN1(n488), .IN2(keyinput51), .Q(n485) );
  NAND2X0 U543 ( .IN1(n489), .IN2(n476), .QN(n488) );
  XNOR2X1 U544 ( .IN1(n490), .IN2(keyinput43), .Q(n476) );
  NAND2X0 U545 ( .IN1(n491), .IN2(n492), .QN(n490) );
  XOR2X1 U546 ( .IN1(keyinput31), .IN2(n493), .Q(n492) );
  AND2X1 U547 ( .IN1(n494), .IN2(n495), .Q(n493) );
  XOR2X1 U548 ( .IN1(n496), .IN2(keyinput30), .Q(n491) );
  NAND2X0 U549 ( .IN1(n495), .IN2(n497), .QN(n496) );
  XOR2X1 U550 ( .IN1(n498), .IN2(keyinput19), .Q(n495) );
  NAND2X0 U551 ( .IN1(n497), .IN2(n494), .QN(n498) );
  XOR3X1 U552 ( .IN1(keyinput7), .IN2(G16), .IN3(G15), .Q(n494) );
  XOR3X1 U553 ( .IN1(keyinput6), .IN2(G14), .IN3(G13), .Q(n497) );
  NOR2X0 U554 ( .IN1(n324), .IN2(n328), .QN(n346) );
  INVX0 U555 ( .INP(n315), .ZN(n328) );
  MUX21X1 U556 ( .IN1(n499), .IN2(n500), .S(n501), .Q(n315) );
  XOR3X1 U557 ( .IN1(G21), .IN2(G17), .IN3(n502), .Q(n501) );
  XNOR2X1 U558 ( .IN1(G29), .IN2(n503), .Q(n502) );
  INVX0 U559 ( .INP(G25), .ZN(n503) );
  XOR2X1 U560 ( .IN1(n504), .IN2(n505), .Q(n500) );
  XNOR2X1 U561 ( .IN1(n504), .IN2(n505), .Q(n499) );
  NAND2X0 U562 ( .IN1(G37), .IN2(G41), .QN(n505) );
  NAND2X0 U563 ( .IN1(n506), .IN2(n507), .QN(n504) );
  XOR2X1 U564 ( .IN1(n508), .IN2(keyinput56), .Q(n507) );
  NAND2X0 U565 ( .IN1(n509), .IN2(n510), .QN(n508) );
  XOR2X1 U566 ( .IN1(n511), .IN2(keyinput57), .Q(n506) );
  NAND2X0 U567 ( .IN1(n509), .IN2(n489), .QN(n511) );
  XOR2X1 U568 ( .IN1(n512), .IN2(keyinput48), .Q(n509) );
  NAND2X0 U569 ( .IN1(n489), .IN2(n510), .QN(n512) );
  INVX0 U570 ( .INP(n487), .ZN(n489) );
  XNOR2X1 U571 ( .IN1(n513), .IN2(keyinput41), .Q(n487) );
  NAND2X0 U572 ( .IN1(n514), .IN2(n515), .QN(n513) );
  XOR2X1 U573 ( .IN1(keyinput27), .IN2(n516), .Q(n515) );
  AND2X1 U574 ( .IN1(n517), .IN2(n518), .Q(n516) );
  XOR2X1 U575 ( .IN1(n519), .IN2(keyinput26), .Q(n514) );
  NAND2X0 U576 ( .IN1(n518), .IN2(n520), .QN(n519) );
  XOR2X1 U577 ( .IN1(n521), .IN2(keyinput17), .Q(n518) );
  NAND2X0 U578 ( .IN1(n517), .IN2(n520), .QN(n521) );
  XOR3X1 U579 ( .IN1(keyinput2), .IN2(G6), .IN3(G5), .Q(n520) );
  XNOR3X1 U580 ( .IN1(keyinput3), .IN2(G8), .IN3(G7), .Q(n517) );
  INVX0 U581 ( .INP(n311), .ZN(n324) );
  MUX21X1 U582 ( .IN1(n522), .IN2(n523), .S(n524), .Q(n311) );
  XOR3X1 U583 ( .IN1(G23), .IN2(G19), .IN3(n525), .Q(n524) );
  XNOR2X1 U584 ( .IN1(G31), .IN2(n526), .Q(n525) );
  INVX0 U585 ( .INP(G27), .ZN(n526) );
  NAND2X0 U586 ( .IN1(n527), .IN2(n528), .QN(n523) );
  AND2X1 U587 ( .IN1(n528), .IN2(n527), .Q(n522) );
  NAND4X0 U588 ( .IN1(G41), .IN2(G39), .IN3(n529), .IN4(n530), .QN(n527) );
  AO22X1 U589 ( .IN1(G41), .IN2(G39), .IN3(n529), .IN4(n530), .Q(n528) );
  NAND2X0 U590 ( .IN1(n474), .IN2(n531), .QN(n530) );
  INVX0 U591 ( .INP(n510), .ZN(n531) );
  INVX0 U592 ( .INP(n477), .ZN(n474) );
  XOR2X1 U593 ( .IN1(n532), .IN2(keyinput50), .Q(n529) );
  NAND2X0 U594 ( .IN1(n510), .IN2(n477), .QN(n532) );
  XNOR2X1 U595 ( .IN1(n533), .IN2(keyinput42), .Q(n477) );
  NAND2X0 U596 ( .IN1(n534), .IN2(n535), .QN(n533) );
  XOR2X1 U597 ( .IN1(keyinput29), .IN2(n536), .Q(n535) );
  AND2X1 U598 ( .IN1(n537), .IN2(n538), .Q(n536) );
  XOR2X1 U599 ( .IN1(n539), .IN2(keyinput28), .Q(n534) );
  NAND2X0 U600 ( .IN1(n540), .IN2(n537), .QN(n539) );
  XNOR2X1 U601 ( .IN1(n541), .IN2(keyinput18), .Q(n537) );
  NAND2X0 U602 ( .IN1(n538), .IN2(n540), .QN(n541) );
  XNOR3X1 U603 ( .IN1(keyinput5), .IN2(G12), .IN3(G11), .Q(n538) );
  XNOR3X1 U604 ( .IN1(keyinput4), .IN2(G9), .IN3(G10), .Q(n540) );
  XNOR2X1 U605 ( .IN1(n542), .IN2(keyinput40), .Q(n510) );
  NAND2X0 U606 ( .IN1(n543), .IN2(n544), .QN(n542) );
  XOR2X1 U607 ( .IN1(keyinput25), .IN2(n545), .Q(n544) );
  AND2X1 U608 ( .IN1(n546), .IN2(n547), .Q(n545) );
  XOR2X1 U609 ( .IN1(n548), .IN2(keyinput24), .Q(n543) );
  NAND2X0 U610 ( .IN1(n547), .IN2(n549), .QN(n548) );
  XOR2X1 U611 ( .IN1(n550), .IN2(keyinput16), .Q(n547) );
  NAND2X0 U612 ( .IN1(n549), .IN2(n546), .QN(n550) );
  XOR3X1 U613 ( .IN1(keyinput1), .IN2(G4), .IN3(G3), .Q(n546) );
  XNOR3X1 U614 ( .IN1(keyinput0), .IN2(G2), .IN3(G1), .Q(n549) );
endmodule

