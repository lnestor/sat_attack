
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572;

  XOR3X1 U344 ( .IN1(keyinput63), .IN2(keyinput60), .IN3(n313), .Q(G1342) );
  NOR2X0 U345 ( .IN1(n314), .IN2(n315), .QN(n313) );
  XOR2X1 U346 ( .IN1(n316), .IN2(keyinput57), .Q(n315) );
  NAND2X0 U347 ( .IN1(n317), .IN2(n318), .QN(n316) );
  XOR2X1 U348 ( .IN1(n319), .IN2(keyinput56), .Q(n314) );
  NAND2X0 U349 ( .IN1(n317), .IN2(G19), .QN(n319) );
  XOR2X1 U350 ( .IN1(n320), .IN2(keyinput51), .Q(n317) );
  NAND2X0 U351 ( .IN1(n318), .IN2(G19), .QN(n320) );
  XOR2X1 U352 ( .IN1(n321), .IN2(keyinput47), .Q(n318) );
  NAND2X0 U353 ( .IN1(n322), .IN2(n323), .QN(n321) );
  XNOR2X1 U354 ( .IN1(G32), .IN2(n324), .Q(G1355) );
  NOR2X0 U355 ( .IN1(n325), .IN2(n326), .QN(n324) );
  XNOR2X1 U356 ( .IN1(G31), .IN2(n327), .Q(G1354) );
  NOR2X0 U357 ( .IN1(n328), .IN2(n326), .QN(n327) );
  XNOR2X1 U358 ( .IN1(G30), .IN2(n329), .Q(G1353) );
  NOR2X0 U359 ( .IN1(n330), .IN2(n326), .QN(n329) );
  XNOR2X1 U360 ( .IN1(G29), .IN2(n331), .Q(G1352) );
  NOR2X0 U361 ( .IN1(n332), .IN2(n326), .QN(n331) );
  NAND4X0 U362 ( .IN1(n333), .IN2(n334), .IN3(n335), .IN4(n336), .QN(n326) );
  XNOR2X1 U363 ( .IN1(G28), .IN2(n337), .Q(G1351) );
  NOR2X0 U364 ( .IN1(n325), .IN2(n338), .QN(n337) );
  XNOR2X1 U365 ( .IN1(G27), .IN2(n339), .Q(G1350) );
  NOR2X0 U366 ( .IN1(n328), .IN2(n338), .QN(n339) );
  XNOR2X1 U367 ( .IN1(G26), .IN2(n340), .Q(G1349) );
  NOR2X0 U368 ( .IN1(n330), .IN2(n338), .QN(n340) );
  XNOR2X1 U369 ( .IN1(G25), .IN2(n341), .Q(G1348) );
  NOR2X0 U370 ( .IN1(n332), .IN2(n338), .QN(n341) );
  NAND4X0 U371 ( .IN1(n342), .IN2(n333), .IN3(n343), .IN4(n344), .QN(n338) );
  NOR2X0 U372 ( .IN1(n345), .IN2(n346), .QN(n343) );
  XNOR2X1 U373 ( .IN1(G24), .IN2(n347), .Q(G1347) );
  NOR2X0 U374 ( .IN1(n325), .IN2(n348), .QN(n347) );
  XNOR2X1 U375 ( .IN1(G23), .IN2(n349), .Q(G1346) );
  NOR2X0 U376 ( .IN1(n328), .IN2(n348), .QN(n349) );
  XNOR2X1 U377 ( .IN1(G22), .IN2(n350), .Q(G1345) );
  NOR2X0 U378 ( .IN1(n330), .IN2(n348), .QN(n350) );
  XNOR2X1 U379 ( .IN1(G21), .IN2(n351), .Q(G1344) );
  NOR2X0 U380 ( .IN1(n332), .IN2(n348), .QN(n351) );
  NAND4X0 U381 ( .IN1(n346), .IN2(n333), .IN3(n352), .IN4(n345), .QN(n348) );
  NOR2X0 U382 ( .IN1(n344), .IN2(n342), .QN(n352) );
  XNOR2X1 U383 ( .IN1(G20), .IN2(n353), .Q(G1343) );
  AND2X1 U384 ( .IN1(n354), .IN2(n323), .Q(n353) );
  XNOR2X1 U385 ( .IN1(G16), .IN2(n355), .Q(G1339) );
  NOR2X0 U386 ( .IN1(n356), .IN2(n357), .QN(n355) );
  XNOR2X1 U387 ( .IN1(G15), .IN2(n358), .Q(G1338) );
  NOR2X0 U388 ( .IN1(n335), .IN2(n357), .QN(n358) );
  XNOR2X1 U389 ( .IN1(G14), .IN2(n359), .Q(G1337) );
  NOR2X0 U390 ( .IN1(n360), .IN2(n357), .QN(n359) );
  XNOR2X1 U391 ( .IN1(G13), .IN2(n361), .Q(G1336) );
  NOR2X0 U392 ( .IN1(n336), .IN2(n357), .QN(n361) );
  NAND3X0 U393 ( .IN1(n354), .IN2(n362), .IN3(n363), .QN(n357) );
  XOR2X1 U394 ( .IN1(n364), .IN2(G12), .Q(G1335) );
  NAND2X0 U395 ( .IN1(n365), .IN2(n346), .QN(n364) );
  XOR2X1 U396 ( .IN1(n366), .IN2(G11), .Q(G1334) );
  NAND2X0 U397 ( .IN1(n365), .IN2(n344), .QN(n366) );
  XOR2X1 U398 ( .IN1(n367), .IN2(G10), .Q(G1333) );
  NAND2X0 U399 ( .IN1(n365), .IN2(n342), .QN(n367) );
  OA22X1 U400 ( .IN1(n368), .IN2(n369), .IN3(n370), .IN4(n369), .Q(G1332) );
  XNOR2X1 U401 ( .IN1(n371), .IN2(keyinput48), .Q(n369) );
  OR2X1 U402 ( .IN1(n368), .IN2(n370), .Q(n371) );
  NAND2X0 U403 ( .IN1(n365), .IN2(n345), .QN(n368) );
  AND3X1 U404 ( .IN1(n372), .IN2(n332), .IN3(n373), .Q(n365) );
  XOR2X1 U405 ( .IN1(n374), .IN2(n375), .Q(G1331) );
  NOR2X0 U406 ( .IN1(n356), .IN2(n376), .QN(n375) );
  XOR2X1 U407 ( .IN1(n377), .IN2(n378), .Q(G1330) );
  NOR2X0 U408 ( .IN1(n335), .IN2(n376), .QN(n378) );
  XOR2X1 U409 ( .IN1(n379), .IN2(n380), .Q(G1329) );
  NOR2X0 U410 ( .IN1(n360), .IN2(n376), .QN(n380) );
  XOR2X1 U411 ( .IN1(n381), .IN2(n382), .Q(G1328) );
  NOR2X0 U412 ( .IN1(n336), .IN2(n376), .QN(n382) );
  NAND4X0 U413 ( .IN1(n383), .IN2(n384), .IN3(n354), .IN4(n362), .QN(n376) );
  XOR2X1 U414 ( .IN1(n385), .IN2(G4), .Q(G1327) );
  NAND2X0 U415 ( .IN1(n386), .IN2(n346), .QN(n385) );
  XOR2X1 U416 ( .IN1(n387), .IN2(G3), .Q(G1326) );
  NAND2X0 U417 ( .IN1(n386), .IN2(n344), .QN(n387) );
  XOR2X1 U418 ( .IN1(n388), .IN2(G2), .Q(G1325) );
  NAND2X0 U419 ( .IN1(n386), .IN2(n342), .QN(n388) );
  XOR2X1 U420 ( .IN1(n389), .IN2(G1), .Q(G1324) );
  NAND2X0 U421 ( .IN1(n386), .IN2(n345), .QN(n389) );
  AND3X1 U422 ( .IN1(n383), .IN2(n330), .IN3(n373), .Q(n386) );
  AND3X1 U423 ( .IN1(n325), .IN2(n362), .IN3(n322), .Q(n373) );
  NAND2X0 U424 ( .IN1(n390), .IN2(n391), .QN(n362) );
  OR3X1 U425 ( .IN1(n342), .IN2(n392), .IN3(n346), .Q(n391) );
  OR3X1 U426 ( .IN1(n345), .IN2(n334), .IN3(n344), .Q(n390) );
  NOR2X0 U427 ( .IN1(n360), .IN2(n356), .QN(n334) );
  XOR3X1 U428 ( .IN1(keyinput62), .IN2(keyinput59), .IN3(n393), .Q(G1341) );
  NAND2X0 U429 ( .IN1(n394), .IN2(n395), .QN(n393) );
  XOR2X1 U430 ( .IN1(n396), .IN2(keyinput54), .Q(n395) );
  NAND2X0 U431 ( .IN1(G18), .IN2(n397), .QN(n396) );
  XOR2X1 U432 ( .IN1(n398), .IN2(keyinput55), .Q(n394) );
  NAND2X0 U433 ( .IN1(n399), .IN2(n397), .QN(n398) );
  XNOR2X1 U434 ( .IN1(n400), .IN2(keyinput50), .Q(n397) );
  NAND2X0 U435 ( .IN1(n399), .IN2(G18), .QN(n400) );
  XOR2X1 U436 ( .IN1(n401), .IN2(keyinput46), .Q(n399) );
  NAND2X0 U437 ( .IN1(n372), .IN2(n323), .QN(n401) );
  XOR3X1 U438 ( .IN1(keyinput61), .IN2(keyinput58), .IN3(n402), .Q(G1340) );
  NOR2X0 U439 ( .IN1(n403), .IN2(n404), .QN(n402) );
  XOR2X1 U440 ( .IN1(keyinput52), .IN2(n405), .Q(n404) );
  AND2X1 U441 ( .IN1(G17), .IN2(n406), .Q(n405) );
  XOR2X1 U442 ( .IN1(n407), .IN2(keyinput53), .Q(n403) );
  NAND2X0 U443 ( .IN1(n406), .IN2(n408), .QN(n407) );
  XOR2X1 U444 ( .IN1(n409), .IN2(keyinput49), .Q(n406) );
  NAND2X0 U445 ( .IN1(n408), .IN2(G17), .QN(n409) );
  XOR2X1 U446 ( .IN1(n410), .IN2(keyinput45), .Q(n408) );
  NAND2X0 U447 ( .IN1(n383), .IN2(n323), .QN(n410) );
  XNOR2X1 U448 ( .IN1(n411), .IN2(keyinput44), .Q(n323) );
  NAND4X0 U449 ( .IN1(n333), .IN2(n392), .IN3(n356), .IN4(n360), .QN(n411) );
  INVX0 U450 ( .INP(n342), .ZN(n360) );
  MUX21X1 U451 ( .IN1(n412), .IN2(n413), .S(n414), .Q(n342) );
  XOR3X1 U452 ( .IN1(G14), .IN2(G10), .IN3(n415), .Q(n414) );
  XOR2X1 U453 ( .IN1(G6), .IN2(G2), .Q(n415) );
  NAND2X0 U454 ( .IN1(n416), .IN2(n417), .QN(n413) );
  AND2X1 U455 ( .IN1(n417), .IN2(n416), .Q(n412) );
  NAND3X0 U456 ( .IN1(G41), .IN2(n418), .IN3(G34), .QN(n416) );
  AO21X1 U457 ( .IN1(G34), .IN2(G41), .IN3(n418), .Q(n417) );
  XOR2X1 U458 ( .IN1(n419), .IN2(n420), .Q(n418) );
  INVX0 U459 ( .INP(n346), .ZN(n356) );
  MUX21X1 U460 ( .IN1(n421), .IN2(n422), .S(n423), .Q(n346) );
  XOR3X1 U461 ( .IN1(G16), .IN2(G12), .IN3(n424), .Q(n423) );
  XOR2X1 U462 ( .IN1(G8), .IN2(G4), .Q(n424) );
  NAND2X0 U463 ( .IN1(n425), .IN2(n426), .QN(n422) );
  AND2X1 U464 ( .IN1(n426), .IN2(n425), .Q(n421) );
  NAND3X0 U465 ( .IN1(G41), .IN2(n427), .IN3(G36), .QN(n425) );
  AO21X1 U466 ( .IN1(G36), .IN2(G41), .IN3(n427), .Q(n426) );
  XOR2X1 U467 ( .IN1(n420), .IN2(n428), .Q(n427) );
  XNOR3X1 U468 ( .IN1(G30), .IN2(G29), .IN3(n429), .Q(n420) );
  XNOR2X1 U469 ( .IN1(G31), .IN2(G32), .Q(n429) );
  NOR2X0 U470 ( .IN1(n336), .IN2(n335), .QN(n392) );
  INVX0 U471 ( .INP(n344), .ZN(n335) );
  MUX21X1 U472 ( .IN1(n430), .IN2(n431), .S(n432), .Q(n344) );
  XOR3X1 U473 ( .IN1(G15), .IN2(G11), .IN3(n433), .Q(n432) );
  XOR2X1 U474 ( .IN1(G7), .IN2(G3), .Q(n433) );
  NAND2X0 U475 ( .IN1(n434), .IN2(n435), .QN(n431) );
  AND2X1 U476 ( .IN1(n435), .IN2(n434), .Q(n430) );
  NAND3X0 U477 ( .IN1(G41), .IN2(n436), .IN3(G35), .QN(n434) );
  AO21X1 U478 ( .IN1(G35), .IN2(G41), .IN3(n436), .Q(n435) );
  XOR2X1 U479 ( .IN1(n419), .IN2(n437), .Q(n436) );
  XNOR3X1 U480 ( .IN1(G26), .IN2(G25), .IN3(n438), .Q(n419) );
  XNOR2X1 U481 ( .IN1(G27), .IN2(G28), .Q(n438) );
  INVX0 U482 ( .INP(n345), .ZN(n336) );
  MUX21X1 U483 ( .IN1(n439), .IN2(n440), .S(n441), .Q(n345) );
  XOR3X1 U484 ( .IN1(G5), .IN2(G1), .IN3(n442), .Q(n441) );
  OA21X1 U485 ( .IN1(G13), .IN2(G9), .IN3(n443), .Q(n442) );
  XOR2X1 U486 ( .IN1(keyinput4), .IN2(n444), .Q(n443) );
  AND2X1 U487 ( .IN1(G9), .IN2(G13), .Q(n444) );
  NAND2X0 U488 ( .IN1(n445), .IN2(n446), .QN(n440) );
  AND2X1 U489 ( .IN1(n446), .IN2(n445), .Q(n439) );
  NAND3X0 U490 ( .IN1(G41), .IN2(n447), .IN3(G33), .QN(n445) );
  AO21X1 U491 ( .IN1(G33), .IN2(G41), .IN3(n447), .Q(n446) );
  XOR2X1 U492 ( .IN1(n428), .IN2(n437), .Q(n447) );
  XNOR3X1 U493 ( .IN1(G18), .IN2(G17), .IN3(n448), .Q(n437) );
  XNOR2X1 U494 ( .IN1(G19), .IN2(G20), .Q(n448) );
  XNOR3X1 U495 ( .IN1(G22), .IN2(G21), .IN3(n449), .Q(n428) );
  XNOR2X1 U496 ( .IN1(G23), .IN2(G24), .Q(n449) );
  XNOR2X1 U497 ( .IN1(keyinput43), .IN2(n450), .Q(n333) );
  NOR3X0 U498 ( .IN1(n451), .IN2(n452), .IN3(n453), .QN(n450) );
  MUX21X1 U499 ( .IN1(n454), .IN2(n455), .S(n332), .Q(n453) );
  NAND3X0 U500 ( .IN1(n456), .IN2(n457), .IN3(n458), .QN(n455) );
  MUX21X1 U501 ( .IN1(n459), .IN2(n460), .S(n330), .Q(n458) );
  NAND3X0 U502 ( .IN1(n322), .IN2(n461), .IN3(n462), .QN(n460) );
  INVX0 U503 ( .INP(keyinput40), .ZN(n461) );
  NAND3X0 U504 ( .IN1(n328), .IN2(n463), .IN3(n464), .QN(n459) );
  INVX0 U505 ( .INP(keyinput41), .ZN(n463) );
  INVX0 U506 ( .INP(n322), .ZN(n328) );
  INVX0 U507 ( .INP(keyinput42), .ZN(n457) );
  NAND2X0 U508 ( .IN1(keyinput39), .IN2(n384), .QN(n456) );
  NOR2X0 U509 ( .IN1(keyinput42), .IN2(n465), .QN(n454) );
  AND2X1 U510 ( .IN1(n465), .IN2(keyinput42), .Q(n452) );
  NAND2X0 U511 ( .IN1(n466), .IN2(n384), .QN(n465) );
  XOR2X1 U512 ( .IN1(n325), .IN2(keyinput38), .Q(n466) );
  AO222X1 U513 ( .IN1(n467), .IN2(n468), .IN3(keyinput41), .IN4(n469), .IN5(
        keyinput40), .IN6(n470), .Q(n451) );
  NAND4X0 U514 ( .IN1(n322), .IN2(n330), .IN3(n332), .IN4(n462), .QN(n470) );
  XOR2X1 U515 ( .IN1(n354), .IN2(keyinput36), .Q(n462) );
  NAND2X0 U516 ( .IN1(n363), .IN2(n464), .QN(n469) );
  XOR2X1 U517 ( .IN1(n354), .IN2(keyinput37), .Q(n464) );
  INVX0 U518 ( .INP(n325), .ZN(n354) );
  XOR2X1 U519 ( .IN1(n471), .IN2(keyinput35), .Q(n325) );
  NAND2X0 U520 ( .IN1(n472), .IN2(n473), .QN(n471) );
  XOR2X1 U521 ( .IN1(n474), .IN2(keyinput33), .Q(n473) );
  NAND2X0 U522 ( .IN1(n475), .IN2(n476), .QN(n474) );
  XOR2X1 U523 ( .IN1(n477), .IN2(keyinput32), .Q(n472) );
  NAND2X0 U524 ( .IN1(n476), .IN2(n478), .QN(n477) );
  XNOR2X1 U525 ( .IN1(n479), .IN2(keyinput31), .Q(n476) );
  NAND2X0 U526 ( .IN1(n475), .IN2(n478), .QN(n479) );
  AO21X1 U527 ( .IN1(n480), .IN2(n481), .IN3(n482), .Q(n478) );
  XOR2X1 U528 ( .IN1(keyinput20), .IN2(n483), .Q(n482) );
  NOR2X0 U529 ( .IN1(n480), .IN2(n481), .QN(n483) );
  XOR2X1 U530 ( .IN1(G28), .IN2(G32), .Q(n481) );
  XNOR2X1 U531 ( .IN1(G20), .IN2(G24), .Q(n480) );
  XOR2X1 U532 ( .IN1(n484), .IN2(keyinput30), .Q(n475) );
  NAND2X0 U533 ( .IN1(n485), .IN2(n486), .QN(n484) );
  XOR2X1 U534 ( .IN1(keyinput28), .IN2(n487), .Q(n486) );
  NOR2X0 U535 ( .IN1(n488), .IN2(n489), .QN(n487) );
  XOR2X1 U536 ( .IN1(keyinput29), .IN2(n490), .Q(n485) );
  NOR2X0 U537 ( .IN1(n488), .IN2(n491), .QN(n490) );
  XNOR2X1 U538 ( .IN1(keyinput26), .IN2(n492), .Q(n491) );
  XOR2X1 U539 ( .IN1(n493), .IN2(keyinput27), .Q(n488) );
  NAND2X0 U540 ( .IN1(n494), .IN2(n495), .QN(n493) );
  XOR2X1 U541 ( .IN1(keyinput26), .IN2(n492), .Q(n495) );
  AND2X1 U542 ( .IN1(n496), .IN2(n497), .Q(n492) );
  XOR2X1 U543 ( .IN1(keyinput24), .IN2(n498), .Q(n497) );
  NOR2X0 U544 ( .IN1(n499), .IN2(n500), .QN(n498) );
  XOR2X1 U545 ( .IN1(keyinput25), .IN2(n501), .Q(n496) );
  NOR2X0 U546 ( .IN1(n502), .IN2(n500), .QN(n501) );
  XNOR2X1 U547 ( .IN1(n503), .IN2(keyinput23), .Q(n500) );
  OR2X1 U548 ( .IN1(n502), .IN2(n499), .Q(n503) );
  INVX0 U549 ( .INP(n489), .ZN(n494) );
  NAND2X0 U550 ( .IN1(G40), .IN2(G41), .QN(n489) );
  NOR3X0 U551 ( .IN1(n322), .IN2(n383), .IN3(n330), .QN(n363) );
  INVX0 U552 ( .INP(n372), .ZN(n330) );
  INVX0 U553 ( .INP(keyinput39), .ZN(n468) );
  NAND2X0 U554 ( .IN1(n384), .IN2(n332), .QN(n467) );
  INVX0 U555 ( .INP(n383), .ZN(n332) );
  NOR2X0 U556 ( .IN1(n322), .IN2(n372), .QN(n384) );
  XOR2X1 U557 ( .IN1(n504), .IN2(n505), .Q(n372) );
  XOR3X1 U558 ( .IN1(G22), .IN2(G18), .IN3(n506), .Q(n505) );
  OA22X1 U559 ( .IN1(n507), .IN2(n508), .IN3(n509), .IN4(n510), .Q(n506) );
  XOR2X1 U560 ( .IN1(n502), .IN2(n511), .Q(n510) );
  AND2X1 U561 ( .IN1(G41), .IN2(G38), .Q(n509) );
  NAND2X0 U562 ( .IN1(G38), .IN2(G41), .QN(n508) );
  XOR2X1 U563 ( .IN1(n502), .IN2(n512), .Q(n507) );
  XNOR2X1 U564 ( .IN1(n513), .IN2(keyinput22), .Q(n502) );
  NAND2X0 U565 ( .IN1(n514), .IN2(n515), .QN(n513) );
  XOR2X1 U566 ( .IN1(n516), .IN2(keyinput19), .Q(n515) );
  NAND2X0 U567 ( .IN1(n517), .IN2(n518), .QN(n516) );
  XOR2X1 U568 ( .IN1(n519), .IN2(keyinput18), .Q(n514) );
  NAND2X0 U569 ( .IN1(n520), .IN2(n517), .QN(n519) );
  XNOR2X1 U570 ( .IN1(n521), .IN2(keyinput15), .Q(n517) );
  NAND2X0 U571 ( .IN1(n520), .IN2(n518), .QN(n521) );
  XNOR2X1 U572 ( .IN1(n522), .IN2(keyinput13), .Q(n518) );
  NAND2X0 U573 ( .IN1(n523), .IN2(n524), .QN(n522) );
  XOR2X1 U574 ( .IN1(keyinput10), .IN2(n525), .Q(n524) );
  AND2X1 U575 ( .IN1(n526), .IN2(G16), .Q(n525) );
  XOR2X1 U576 ( .IN1(n527), .IN2(keyinput9), .Q(n523) );
  NAND2X0 U577 ( .IN1(G15), .IN2(n526), .QN(n527) );
  XNOR2X1 U578 ( .IN1(n528), .IN2(keyinput3), .Q(n526) );
  NAND2X0 U579 ( .IN1(G16), .IN2(G15), .QN(n528) );
  XOR2X1 U580 ( .IN1(n529), .IN2(keyinput12), .Q(n520) );
  NAND2X0 U581 ( .IN1(n530), .IN2(n531), .QN(n529) );
  XOR2X1 U582 ( .IN1(keyinput8), .IN2(n532), .Q(n531) );
  AND2X1 U583 ( .IN1(n533), .IN2(G14), .Q(n532) );
  XOR2X1 U584 ( .IN1(n534), .IN2(keyinput7), .Q(n530) );
  NAND2X0 U585 ( .IN1(G13), .IN2(n533), .QN(n534) );
  XNOR2X1 U586 ( .IN1(n535), .IN2(keyinput2), .Q(n533) );
  NAND2X0 U587 ( .IN1(G14), .IN2(G13), .QN(n535) );
  XNOR3X1 U588 ( .IN1(keyinput34), .IN2(G30), .IN3(G26), .Q(n504) );
  MUX21X1 U589 ( .IN1(n536), .IN2(n537), .S(n538), .Q(n322) );
  XOR3X1 U590 ( .IN1(G23), .IN2(G19), .IN3(n539), .Q(n538) );
  XOR2X1 U591 ( .IN1(G31), .IN2(G27), .Q(n539) );
  NAND2X0 U592 ( .IN1(n540), .IN2(n541), .QN(n537) );
  AND2X1 U593 ( .IN1(n541), .IN2(n540), .Q(n536) );
  NAND3X0 U594 ( .IN1(G39), .IN2(n542), .IN3(G41), .QN(n540) );
  AO21X1 U595 ( .IN1(G41), .IN2(G39), .IN3(n542), .Q(n541) );
  XOR2X1 U596 ( .IN1(n543), .IN2(n512), .Q(n542) );
  INVX0 U597 ( .INP(n511), .ZN(n512) );
  XOR3X1 U598 ( .IN1(G11), .IN2(G10), .IN3(n544), .Q(n511) );
  XOR2X1 U599 ( .IN1(G12), .IN2(n370), .Q(n544) );
  INVX0 U600 ( .INP(G9), .ZN(n370) );
  MUX21X1 U601 ( .IN1(n545), .IN2(n546), .S(n547), .Q(n383) );
  XOR3X1 U602 ( .IN1(G21), .IN2(G17), .IN3(n548), .Q(n547) );
  XOR2X1 U603 ( .IN1(G29), .IN2(G25), .Q(n548) );
  NAND2X0 U604 ( .IN1(n549), .IN2(n550), .QN(n546) );
  AND2X1 U605 ( .IN1(n550), .IN2(n549), .Q(n545) );
  NAND3X0 U606 ( .IN1(G37), .IN2(G41), .IN3(n551), .QN(n549) );
  AO21X1 U607 ( .IN1(G37), .IN2(G41), .IN3(n551), .Q(n550) );
  XNOR2X1 U608 ( .IN1(n499), .IN2(n543), .Q(n551) );
  XNOR3X1 U609 ( .IN1(G2), .IN2(G1), .IN3(n552), .Q(n543) );
  XNOR2X1 U610 ( .IN1(G3), .IN2(G4), .Q(n552) );
  XNOR2X1 U611 ( .IN1(n553), .IN2(keyinput21), .Q(n499) );
  NAND2X0 U612 ( .IN1(n554), .IN2(n555), .QN(n553) );
  XOR2X1 U613 ( .IN1(keyinput16), .IN2(n556), .Q(n555) );
  NOR2X0 U614 ( .IN1(n557), .IN2(n558), .QN(n556) );
  XNOR2X1 U615 ( .IN1(keyinput11), .IN2(n559), .Q(n558) );
  XOR2X1 U616 ( .IN1(n560), .IN2(keyinput17), .Q(n554) );
  NAND2X0 U617 ( .IN1(n561), .IN2(n562), .QN(n560) );
  INVX0 U618 ( .INP(n557), .ZN(n562) );
  XOR2X1 U619 ( .IN1(n563), .IN2(keyinput14), .Q(n557) );
  NAND2X0 U620 ( .IN1(n564), .IN2(n561), .QN(n563) );
  XOR2X1 U621 ( .IN1(n559), .IN2(keyinput11), .Q(n564) );
  NAND2X0 U622 ( .IN1(n565), .IN2(n566), .QN(n559) );
  XOR2X1 U623 ( .IN1(keyinput5), .IN2(n567), .Q(n566) );
  NOR2X0 U624 ( .IN1(n568), .IN2(n381), .QN(n567) );
  INVX0 U625 ( .INP(G5), .ZN(n381) );
  XOR2X1 U626 ( .IN1(keyinput6), .IN2(n569), .Q(n565) );
  NOR2X0 U627 ( .IN1(n568), .IN2(n379), .QN(n569) );
  INVX0 U628 ( .INP(G6), .ZN(n379) );
  XOR2X1 U629 ( .IN1(n570), .IN2(keyinput0), .Q(n568) );
  NAND2X0 U630 ( .IN1(G6), .IN2(G5), .QN(n570) );
  AOI21X1 U631 ( .IN1(n377), .IN2(n374), .IN3(n571), .QN(n561) );
  XOR2X1 U632 ( .IN1(keyinput1), .IN2(n572), .Q(n571) );
  NOR2X0 U633 ( .IN1(n377), .IN2(n374), .QN(n572) );
  INVX0 U634 ( .INP(G8), .ZN(n374) );
  INVX0 U635 ( .INP(G7), .ZN(n377) );
endmodule

