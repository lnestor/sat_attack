
module c1908 ( N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, 
        N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, 
        N85, N88, N91, N94, N99, N104, N2753, N2754, N2755, N2756, N2762, 
        N2767, N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, 
        N2787, N2811, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31 );
  input N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43,
         N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88,
         N91, N94, N99, N104, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31;
  output N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781,
         N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888,
         N2889, N2890, N2891, N2892, N2899;
  wire   n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435;

  NOR2X0 U252 ( .IN1(n244), .IN2(n245), .QN(N2899) );
  XOR3X1 U253 ( .IN1(n246), .IN2(n247), .IN3(n248), .Q(n245) );
  NAND2X0 U254 ( .IN1(n249), .IN2(N79), .QN(n247) );
  XOR3X1 U255 ( .IN1(n250), .IN2(n251), .IN3(n252), .Q(N2892) );
  NAND2X0 U256 ( .IN1(n253), .IN2(n254), .QN(n252) );
  OA21X1 U257 ( .IN1(N66), .IN2(n254), .IN3(n255), .Q(n251) );
  NOR2X0 U258 ( .IN1(n256), .IN2(n257), .QN(n250) );
  XOR2X1 U259 ( .IN1(n258), .IN2(n259), .Q(n257) );
  INVX0 U260 ( .INP(n255), .ZN(n256) );
  NAND2X0 U261 ( .IN1(N104), .IN2(n260), .QN(n255) );
  XOR3X1 U262 ( .IN1(n261), .IN2(n262), .IN3(n263), .Q(N2891) );
  AND2X1 U263 ( .IN1(n254), .IN2(n264), .Q(n263) );
  AOI21X1 U264 ( .IN1(N63), .IN2(N88), .IN3(n254), .QN(n262) );
  OA21X1 U265 ( .IN1(n254), .IN2(n265), .IN3(n266), .Q(n261) );
  XOR2X1 U266 ( .IN1(keyinput1), .IN2(N88), .Q(n265) );
  NOR2X0 U267 ( .IN1(n244), .IN2(n267), .QN(N2890) );
  XNOR2X1 U268 ( .IN1(n268), .IN2(n269), .Q(n267) );
  NAND2X0 U269 ( .IN1(n249), .IN2(n270), .QN(n268) );
  NOR2X0 U270 ( .IN1(n244), .IN2(n271), .QN(N2889) );
  XOR3X1 U271 ( .IN1(keyinput31), .IN2(n272), .IN3(n273), .Q(n271) );
  NAND2X0 U272 ( .IN1(N85), .IN2(n249), .QN(n272) );
  NOR2X0 U273 ( .IN1(n244), .IN2(n274), .QN(N2888) );
  XOR2X1 U274 ( .IN1(n275), .IN2(n276), .Q(n274) );
  NAND3X0 U275 ( .IN1(n249), .IN2(N82), .IN3(keyinput13), .QN(n276) );
  NOR2X0 U276 ( .IN1(n244), .IN2(n277), .QN(N2887) );
  XOR2X1 U277 ( .IN1(n278), .IN2(n279), .Q(n277) );
  NAND2X0 U278 ( .IN1(n249), .IN2(N76), .QN(n278) );
  NOR2X0 U279 ( .IN1(n244), .IN2(n280), .QN(N2886) );
  XOR3X1 U280 ( .IN1(n281), .IN2(n282), .IN3(n283), .Q(n280) );
  XOR2X1 U281 ( .IN1(n284), .IN2(n285), .Q(n283) );
  NOR2X0 U282 ( .IN1(keyinput15), .IN2(n266), .QN(n285) );
  NAND2X0 U283 ( .IN1(n249), .IN2(n286), .QN(n284) );
  NOR2X0 U284 ( .IN1(n287), .IN2(n288), .QN(n249) );
  OA21X1 U285 ( .IN1(n289), .IN2(n290), .IN3(n291), .Q(n281) );
  XOR2X1 U286 ( .IN1(n292), .IN2(keyinput10), .Q(n291) );
  NOR2X0 U287 ( .IN1(n254), .IN2(N99), .QN(n244) );
  OR2X1 U288 ( .IN1(n293), .IN2(n294), .Q(N2811) );
  NOR4X0 U289 ( .IN1(n295), .IN2(n296), .IN3(n297), .IN4(n298), .QN(n294) );
  INVX0 U290 ( .INP(n299), .ZN(n297) );
  XNOR2X1 U291 ( .IN1(N85), .IN2(n300), .Q(n296) );
  NAND4X0 U292 ( .IN1(n301), .IN2(n302), .IN3(n303), .IN4(n304), .QN(n295) );
  XOR2X1 U293 ( .IN1(keyinput17), .IN2(n305), .Q(n303) );
  XOR2X1 U294 ( .IN1(keyinput16), .IN2(n306), .Q(n302) );
  OA22X1 U295 ( .IN1(N104), .IN2(n307), .IN3(N104), .IN4(N99), .Q(n293) );
  XOR2X1 U296 ( .IN1(n308), .IN2(keyinput30), .Q(n307) );
  NAND2X0 U297 ( .IN1(n288), .IN2(n309), .QN(n308) );
  XNOR2X1 U298 ( .IN1(n310), .IN2(keyinput24), .Q(n309) );
  NAND2X0 U299 ( .IN1(n311), .IN2(n312), .QN(n310) );
  NAND4X0 U300 ( .IN1(n313), .IN2(n314), .IN3(n315), .IN4(n316), .QN(n312) );
  AO221X1 U301 ( .IN1(n317), .IN2(n318), .IN3(n319), .IN4(n299), .IN5(n320), 
        .Q(n316) );
  AO22X1 U302 ( .IN1(n321), .IN2(n299), .IN3(n322), .IN4(n323), .Q(n320) );
  NOR2X0 U303 ( .IN1(n324), .IN2(n325), .QN(n322) );
  INVX0 U304 ( .INP(n318), .ZN(n324) );
  NAND4X0 U305 ( .IN1(n313), .IN2(n318), .IN3(n299), .IN4(n326), .QN(n311) );
  AO222X1 U306 ( .IN1(n315), .IN2(n327), .IN3(n314), .IN4(n328), .IN5(n329), 
        .IN6(n330), .Q(n326) );
  MUX21X1 U307 ( .IN1(n331), .IN2(n315), .S(n332), .Q(n329) );
  NOR2X0 U308 ( .IN1(n264), .IN2(n253), .QN(n288) );
  NAND4X0 U309 ( .IN1(n333), .IN2(n334), .IN3(n335), .IN4(n336), .QN(n253) );
  NOR4X0 U310 ( .IN1(n337), .IN2(n338), .IN3(n339), .IN4(n340), .QN(n336) );
  NOR2X0 U311 ( .IN1(n341), .IN2(n342), .QN(n335) );
  INVX0 U312 ( .INP(n343), .ZN(n341) );
  NAND4X0 U313 ( .IN1(n344), .IN2(n345), .IN3(n346), .IN4(n347), .QN(n264) );
  NOR4X0 U314 ( .IN1(n348), .IN2(n349), .IN3(n350), .IN4(n351), .QN(n347) );
  AND2X1 U315 ( .IN1(n352), .IN2(n353), .Q(n346) );
  XOR2X1 U316 ( .IN1(keyinput22), .IN2(n354), .Q(n344) );
  XOR2X1 U317 ( .IN1(n355), .IN2(n333), .Q(N2787) );
  NAND3X0 U318 ( .IN1(n331), .IN2(n319), .IN3(n356), .QN(n333) );
  XNOR2X1 U319 ( .IN1(N37), .IN2(n334), .Q(N2786) );
  NAND4X0 U320 ( .IN1(n356), .IN2(n318), .IN3(n298), .IN4(n306), .QN(n334) );
  XOR3X1 U321 ( .IN1(keyinput29), .IN2(n342), .IN3(n357), .Q(N2785) );
  NAND2X0 U322 ( .IN1(keyinput27), .IN2(N34), .QN(n357) );
  AND3X1 U323 ( .IN1(n321), .IN2(n328), .IN3(n356), .Q(n342) );
  XOR2X1 U324 ( .IN1(N31), .IN2(n338), .Q(N2784) );
  AND3X1 U325 ( .IN1(n328), .IN2(n319), .IN3(n356), .Q(n338) );
  AND2X1 U326 ( .IN1(n314), .IN2(n358), .Q(n356) );
  AND2X1 U327 ( .IN1(n330), .IN2(n304), .Q(n314) );
  XOR2X1 U328 ( .IN1(n290), .IN2(n343), .Q(N2783) );
  NAND4X0 U329 ( .IN1(n327), .IN2(n359), .IN3(n299), .IN4(n360), .QN(n343) );
  AND2X1 U330 ( .IN1(n319), .IN2(n331), .Q(n360) );
  XNOR2X1 U331 ( .IN1(N22), .IN2(n345), .Q(N2782) );
  NAND4X0 U332 ( .IN1(n361), .IN2(n315), .IN3(n362), .IN4(n305), .QN(n345) );
  XOR2X1 U333 ( .IN1(N19), .IN2(n349), .Q(N2781) );
  AND4X1 U334 ( .IN1(n318), .IN2(n362), .IN3(n298), .IN4(n306), .Q(n349) );
  XOR3X1 U335 ( .IN1(keyinput28), .IN2(N16), .IN3(n363), .Q(N2780) );
  NOR2X0 U336 ( .IN1(keyinput2), .IN2(n364), .QN(n363) );
  XOR2X1 U337 ( .IN1(keyinput23), .IN2(n354), .Q(n364) );
  AND3X1 U338 ( .IN1(n328), .IN2(n362), .IN3(n321), .Q(n354) );
  XOR2X1 U339 ( .IN1(n348), .IN2(n365), .Q(N2779) );
  NOR2X0 U340 ( .IN1(keyinput26), .IN2(n366), .QN(n365) );
  AND3X1 U341 ( .IN1(n319), .IN2(n362), .IN3(n328), .Q(n348) );
  AND2X1 U342 ( .IN1(n367), .IN2(n299), .Q(n362) );
  NOR2X0 U343 ( .IN1(n325), .IN2(n323), .QN(n299) );
  INVX0 U344 ( .INP(n368), .ZN(n323) );
  XNOR3X1 U345 ( .IN1(keyinput21), .IN2(n340), .IN3(N46), .Q(N2768) );
  AND2X1 U346 ( .IN1(n369), .IN2(n319), .Q(n340) );
  XOR2X1 U347 ( .IN1(N43), .IN2(n339), .Q(N2767) );
  AND4X1 U348 ( .IN1(n327), .IN2(n305), .IN3(n328), .IN4(n370), .Q(n339) );
  NOR2X0 U349 ( .IN1(n371), .IN2(n372), .QN(n370) );
  XOR2X1 U350 ( .IN1(N28), .IN2(n337), .Q(N2762) );
  AND2X1 U351 ( .IN1(n369), .IN2(n321), .Q(n337) );
  AND4X1 U352 ( .IN1(n358), .IN2(n327), .IN3(n298), .IN4(n306), .Q(n369) );
  INVX0 U353 ( .INP(n371), .ZN(n358) );
  NAND2X0 U354 ( .IN1(n317), .IN2(n359), .QN(n371) );
  AO21X1 U355 ( .IN1(n373), .IN2(n260), .IN3(n313), .Q(n359) );
  INVX0 U356 ( .INP(N91), .ZN(n260) );
  XNOR2X1 U357 ( .IN1(N10), .IN2(n353), .Q(N2756) );
  NAND3X0 U358 ( .IN1(n374), .IN2(n318), .IN3(n331), .QN(n353) );
  XOR2X1 U359 ( .IN1(n375), .IN2(keyinput20), .Q(n331) );
  NAND2X0 U360 ( .IN1(n376), .IN2(n306), .QN(n375) );
  XNOR2X1 U361 ( .IN1(N7), .IN2(n352), .Q(N2755) );
  NAND3X0 U362 ( .IN1(n315), .IN2(n374), .IN3(n321), .QN(n352) );
  NOR2X0 U363 ( .IN1(n372), .IN2(n305), .QN(n321) );
  AO21X1 U364 ( .IN1(n351), .IN2(n377), .IN3(n378), .Q(N2754) );
  XOR2X1 U365 ( .IN1(keyinput25), .IN2(n379), .Q(n378) );
  NOR2X0 U366 ( .IN1(n351), .IN2(n377), .QN(n379) );
  AND3X1 U367 ( .IN1(n374), .IN2(n319), .IN3(n315), .Q(n351) );
  NOR2X0 U368 ( .IN1(n298), .IN2(n306), .QN(n315) );
  INVX0 U369 ( .INP(n376), .ZN(n298) );
  AND2X1 U370 ( .IN1(n372), .IN2(n305), .Q(n319) );
  INVX0 U371 ( .INP(n361), .ZN(n372) );
  XOR2X1 U372 ( .IN1(N1), .IN2(n350), .Q(N2753) );
  AND3X1 U373 ( .IN1(n318), .IN2(n328), .IN3(n374), .Q(n350) );
  AND2X1 U374 ( .IN1(n317), .IN2(n367), .Q(n374) );
  AND2X1 U375 ( .IN1(n327), .IN2(n380), .Q(n367) );
  AO21X1 U376 ( .IN1(n381), .IN2(n373), .IN3(n313), .Q(n380) );
  OA21X1 U377 ( .IN1(n382), .IN2(n383), .IN3(N99), .Q(n313) );
  NOR2X0 U378 ( .IN1(N104), .IN2(N69), .QN(n383) );
  AND3X1 U379 ( .IN1(N104), .IN2(n384), .IN3(N94), .Q(n373) );
  NAND2X0 U380 ( .IN1(N72), .IN2(N69), .QN(n384) );
  XNOR2X1 U381 ( .IN1(N88), .IN2(keyinput1), .Q(n381) );
  NOR2X0 U382 ( .IN1(n330), .IN2(n332), .QN(n327) );
  INVX0 U383 ( .INP(n304), .ZN(n332) );
  NAND2X0 U384 ( .IN1(N53), .IN2(n385), .QN(n304) );
  XOR2X1 U385 ( .IN1(n301), .IN2(keyinput19), .Q(n330) );
  XOR3X1 U386 ( .IN1(keyinput18), .IN2(n286), .IN3(n386), .Q(n301) );
  NAND2X0 U387 ( .IN1(n387), .IN2(n287), .QN(n386) );
  XNOR3X1 U388 ( .IN1(n282), .IN2(n388), .IN3(n266), .Q(n387) );
  XOR3X1 U389 ( .IN1(n389), .IN2(n390), .IN3(n391), .Q(n266) );
  XNOR3X1 U390 ( .IN1(N22), .IN2(n392), .IN3(N10), .Q(n391) );
  NOR2X0 U391 ( .IN1(keyinput3), .IN2(n393), .QN(n392) );
  OA22X1 U392 ( .IN1(n394), .IN2(n395), .IN3(N1), .IN4(n396), .Q(n389) );
  NOR2X0 U393 ( .IN1(n397), .IN2(n398), .QN(n396) );
  OR2X1 U394 ( .IN1(n399), .IN2(n397), .Q(n395) );
  OA21X1 U395 ( .IN1(n289), .IN2(n400), .IN3(n292), .Q(n388) );
  NAND2X0 U396 ( .IN1(n289), .IN2(n290), .QN(n292) );
  XOR2X1 U397 ( .IN1(keyinput6), .IN2(N25), .Q(n400) );
  NAND2X0 U398 ( .IN1(N63), .IN2(n254), .QN(n282) );
  AND2X1 U399 ( .IN1(N49), .IN2(n385), .Q(n286) );
  OR2X1 U400 ( .IN1(N94), .IN2(N72), .Q(n385) );
  AND2X1 U401 ( .IN1(n325), .IN2(n368), .Q(n317) );
  NAND2X0 U402 ( .IN1(N60), .IN2(n401), .QN(n368) );
  XNOR2X1 U403 ( .IN1(n402), .IN2(N76), .Q(n325) );
  NAND2X0 U404 ( .IN1(n403), .IN2(n287), .QN(n402) );
  XOR2X1 U405 ( .IN1(n279), .IN2(keyinput9), .Q(n403) );
  XOR3X1 U406 ( .IN1(n404), .IN2(n258), .IN3(n405), .Q(n279) );
  XOR3X1 U407 ( .IN1(N40), .IN2(N10), .IN3(n406), .Q(n405) );
  NAND2X0 U408 ( .IN1(N66), .IN2(n254), .QN(n406) );
  OA22X1 U409 ( .IN1(n407), .IN2(n408), .IN3(N1), .IN4(n409), .Q(n404) );
  NOR2X0 U410 ( .IN1(n398), .IN2(n407), .QN(n409) );
  INVX0 U411 ( .INP(n394), .ZN(n398) );
  OR2X1 U412 ( .IN1(n394), .IN2(n399), .Q(n408) );
  NOR2X0 U413 ( .IN1(N1), .IN2(n399), .QN(n394) );
  AND2X1 U414 ( .IN1(N7), .IN2(n377), .Q(n399) );
  MUX21X1 U415 ( .IN1(n397), .IN2(n377), .S(keyinput5), .Q(n407) );
  NOR2X0 U416 ( .IN1(n377), .IN2(N7), .QN(n397) );
  INVX0 U417 ( .INP(N4), .ZN(n377) );
  NOR2X0 U418 ( .IN1(n306), .IN2(n376), .QN(n328) );
  XOR2X1 U419 ( .IN1(n410), .IN2(N79), .Q(n376) );
  NAND2X0 U420 ( .IN1(n411), .IN2(n287), .QN(n410) );
  XOR2X1 U421 ( .IN1(n412), .IN2(n413), .Q(n411) );
  INVX0 U422 ( .INP(n248), .ZN(n413) );
  XOR2X1 U423 ( .IN1(n414), .IN2(N1), .Q(n248) );
  NAND2X0 U424 ( .IN1(N49), .IN2(n382), .QN(n414) );
  NOR2X0 U425 ( .IN1(keyinput7), .IN2(n246), .QN(n412) );
  XNOR3X1 U426 ( .IN1(n390), .IN2(n393), .IN3(n258), .Q(n246) );
  XOR3X1 U427 ( .IN1(N31), .IN2(n415), .IN3(n289), .Q(n258) );
  XOR2X1 U428 ( .IN1(N46), .IN2(n416), .Q(n289) );
  XOR2X1 U429 ( .IN1(N37), .IN2(N34), .Q(n415) );
  XOR2X1 U430 ( .IN1(N13), .IN2(N19), .Q(n390) );
  XOR2X1 U431 ( .IN1(n270), .IN2(n417), .Q(n306) );
  NOR2X0 U432 ( .IN1(N94), .IN2(n269), .QN(n417) );
  XNOR2X1 U433 ( .IN1(n418), .IN2(n419), .Q(n269) );
  XOR3X1 U434 ( .IN1(n420), .IN2(n421), .IN3(n422), .Q(n419) );
  NAND3X0 U435 ( .IN1(N69), .IN2(n254), .IN3(N60), .QN(n422) );
  NAND2X0 U436 ( .IN1(keyinput4), .IN2(n355), .QN(n421) );
  XOR2X1 U437 ( .IN1(N19), .IN2(N10), .Q(n420) );
  XOR3X1 U438 ( .IN1(N28), .IN2(N25), .IN3(n423), .Q(n418) );
  XNOR2X1 U439 ( .IN1(N37), .IN2(N46), .Q(n423) );
  AND2X1 U440 ( .IN1(N56), .IN2(n401), .Q(n270) );
  NAND2X0 U441 ( .IN1(N69), .IN2(n287), .QN(n401) );
  NOR2X0 U442 ( .IN1(n305), .IN2(n361), .QN(n318) );
  XOR2X1 U443 ( .IN1(n300), .IN2(n424), .Q(n361) );
  NOR2X0 U444 ( .IN1(N85), .IN2(keyinput14), .QN(n424) );
  NAND2X0 U445 ( .IN1(n273), .IN2(n287), .QN(n300) );
  XNOR3X1 U446 ( .IN1(n416), .IN2(n425), .IN3(n426), .Q(n273) );
  XOR3X1 U447 ( .IN1(keyinput12), .IN2(N34), .IN3(n427), .Q(n426) );
  NAND2X0 U448 ( .IN1(keyinput8), .IN2(n428), .QN(n427) );
  XNOR3X1 U449 ( .IN1(N7), .IN2(N22), .IN3(n393), .Q(n428) );
  XNOR2X1 U450 ( .IN1(N16), .IN2(keyinput0), .Q(n393) );
  NAND3X0 U451 ( .IN1(N69), .IN2(n254), .IN3(N56), .QN(n425) );
  INVX0 U452 ( .INP(N104), .ZN(n254) );
  XOR2X1 U453 ( .IN1(N28), .IN2(N43), .Q(n416) );
  XNOR2X1 U454 ( .IN1(n429), .IN2(N82), .Q(n305) );
  NAND2X0 U455 ( .IN1(n287), .IN2(n275), .QN(n429) );
  AO21X1 U456 ( .IN1(n430), .IN2(n431), .IN3(n432), .Q(n275) );
  XOR2X1 U457 ( .IN1(keyinput11), .IN2(n433), .Q(n432) );
  NOR2X0 U458 ( .IN1(n430), .IN2(n431), .QN(n433) );
  XOR3X1 U459 ( .IN1(n259), .IN2(n434), .IN3(n435), .Q(n431) );
  XNOR3X1 U460 ( .IN1(N46), .IN2(N43), .IN3(N31), .Q(n435) );
  NAND2X0 U461 ( .IN1(N53), .IN2(n382), .QN(n434) );
  NOR2X0 U462 ( .IN1(N104), .IN2(N72), .QN(n382) );
  XOR2X1 U463 ( .IN1(n355), .IN2(n290), .Q(n259) );
  INVX0 U464 ( .INP(N25), .ZN(n290) );
  INVX0 U465 ( .INP(N40), .ZN(n355) );
  XOR3X1 U466 ( .IN1(N4), .IN2(N22), .IN3(n366), .Q(n430) );
  INVX0 U467 ( .INP(N13), .ZN(n366) );
  INVX0 U468 ( .INP(N94), .ZN(n287) );
endmodule

