// Verilog File 
module c1908_xor_256bit.bench (G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,
keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,
keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,
keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,
keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,
keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,
keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,
keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,
keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,
keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,
keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205,
keyinput206,keyinput207,keyinput208,keyinput209,keyinput210,keyinput211,keyinput212,keyinput213,keyinput214,keyinput215,
keyinput216,keyinput217,keyinput218,keyinput219,keyinput220,keyinput221,keyinput222,keyinput223,keyinput224,keyinput225,
keyinput226,keyinput227,keyinput228,keyinput229,keyinput230,keyinput231,keyinput232,keyinput233,keyinput234,keyinput235,
keyinput236,keyinput237,keyinput238,keyinput239,keyinput240,keyinput241,keyinput242,keyinput243,keyinput244,keyinput245,
keyinput246,keyinput247,keyinput248,keyinput249,keyinput250,keyinput251,keyinput252,keyinput253,keyinput254,keyinput255,
G3,G6,G9,G12,G30,G45,G48,G15,G18,G21,
G24,G27,G33,G36,G39,G42,G75,G51,G54,G60,
G63,G66,G69,G72,G57);

input G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,
keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,
keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,
keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,
keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,
keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,
keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,
keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,
keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,
keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,
keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205,
keyinput206,keyinput207,keyinput208,keyinput209,keyinput210,keyinput211,keyinput212,keyinput213,keyinput214,keyinput215,
keyinput216,keyinput217,keyinput218,keyinput219,keyinput220,keyinput221,keyinput222,keyinput223,keyinput224,keyinput225,
keyinput226,keyinput227,keyinput228,keyinput229,keyinput230,keyinput231,keyinput232,keyinput233,keyinput234,keyinput235,
keyinput236,keyinput237,keyinput238,keyinput239,keyinput240,keyinput241,keyinput242,keyinput243,keyinput244,keyinput245,
keyinput246,keyinput247,keyinput248,keyinput249,keyinput250,keyinput251,keyinput252,keyinput253,keyinput254,keyinput255;


output G3, G6, G9, G12, G30, G45, G48, G15, G18, 
G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, 
G60, G63, G66, G69, G72, G57;

wire G149, G153, G156, G160, G165, G168, G171, G175, G179, 
G184, G188, G191, G194, G198, G202, G206, G231, G233, G241, 
G244, G245, G248, G517, G529, G541, G553, G859, G862, G907, 
G909, G911, G918, G919, G922, G926, G930, G932, G934, G938, 
G943, G947, G949, G1506, G1514, G1522, G1530, G1538, G1546, G1554, 
G1562, G1570, G1578, G1586, G1594, G1602, G1610, G1618, G1626, G1512, 
G1520, G1528, G1536, G1544, xenc200, G1552, xenc231, G1560, xenc33, G1568, 
xenc14, G1576, G1584, xenc5, G1592, G1600, xenc9, G1608, G1616, xenc122, 
G1624, G1632, xenc95, G50, G52, G56, G58, G62, G64, xenc169, 
G251, xenc100, G254, xenc124, G288, G291, G299, G302, xenc0, G318, 
G321, G327, G330, G352, xenc244, G355, G369, xenc145, G382, G385, 
xenc254, G853, G856, xenc176, G893, xenc130, G954, G955, xenc246, G1050, 
G1053, G1176, G1179, G1197, G1207, G1222, G1244, G1278, G1290, G1300, 
G1312, G1332, G1335, G1442, G1450, G1458, G1466, G1474, G1482, xenc15, 
G1490, G1498, G1634, G1644, G1657, G1665, xenc61, G1697, G1705, G1713, 
G1721, G1745, G1753, G1785, G1793, G1814, G1817, G1830, G1833, G1841, 
G1849, G1854, G1857, G1870, G1873, G1878, G1881, G1642, G1652, G1056, 
G1057, G1182, xenc60, G1183, G1211, xenc91, G1298, G1320, xenc111, G1338, 
G1339, xenc141, G457, xenc172, G459, G482, G487, G492, G505, G1456, 
G1448, xenc224, G1472, G1464, G1488, xenc203, G1480, G1504, G1496, xenc184, 
G956, G967, xenc212, G978, G979, G980, G1661, G990, G1669, G1030, 
xenc144, G1701, G1040, xenc152, G1709, G1058, G1717, G1068, G1725, xenc197, 
G1078, G1090, G1100, G1749, G1112, xenc59, G1757, G1154, xenc223, G1789, 
G1166, G1797, xenc67, G1194, G1201, G1204, xenc36, G1820, G1821, xenc229, 
G1230, xenc94, G1836, G1837, G1252, G1256, G1845, G1268, G1853, xenc239, 
G1860, G1861, G1286, G1876, G1877, G1308, xenc44, G1884, G1885, xenc12, 
G1654, G1662, G1694, G1702, xenc29, G1710, G1718, G1726, G1734, G1742, 
G1750, G1782, G1790, G1838, G1846, xenc250, G297, xenc3, G298, G361, 
xenc206, G362, xenc162, G404, G405, G1225, G1226, G1247, xenc165, G1248, 
G1281, G1282, xenc190, G1303, G1304, G1315, xenc154, G1316, xenc155, G998, 
G988, G268, G1038, G1048, G1076, G1066, G1098, xenc195, G1120, G1174, 
G363, G1210, G373, G1276, xenc161, G406, G565, G566, G614, G615, 
G958, G969, xenc147, G1660, xenc255, G984, G1668, G994, G1700, xenc191, 
G1034, G1708, xenc138, G1044, xenc27, G1716, G1062, G1724, G1072, G1732, 
xenc121, G1086, G1740, xenc53, G1748, xenc177, G1104, xenc25, G1108, G1756, 
xenc96, G1116, G1788, G1158, G1162, G1796, G1170, G1200, G1203, G1227, 
G1249, G1844, G1260, G1264, G1852, G1272, xenc113, G1283, xenc20, xenc69, 
G1305, G1317, G1410, G1418, xenc17, G1426, G1434, xenc222, G269, xenc185, 
G372, xenc205, G983, G993, G1033, G1043, G1061, G1071, G1103, G1115, 
xenc237, G1157, G1169, xenc101, G1184, G1202, G1259, G1271, G1322, xenc248, 
G374, xenc230, xenc102, G396, G1321, G1424, G1416, G1440, G1432, xenc242, 
G985, G995, G1035, G1045, xenc175, G1063, G1073, xenc23, G1105, xenc50, 
G1117, G1159, G1171, G1212, G1231, G1232, G1253, xenc236, G1254, G1261, 
xenc64, xenc109, G1273, G1287, G1288, G1309, G1310, G1192, G397, G1330, 
G1000, G1010, G1233, G1255, xenc18, G1289, xenc136, G1311, G1381, G257, 
G999, G260, G989, G272, G1039, G294, G1049, G305, G1077, xenc128, 
G308, G1067, xenc22, xenc42, G333, G1121, G358, G1175, xenc143, G1220, 
xenc66, xenc123, G388, G1277, G398, xenc215, G1109, G1110, xenc30, G1163, 
G1164, G1234, G1265, G1266, G1822, G1862, xenc115, G1865, xenc92, G258, 
xenc81, G261, G273, xenc13, G1018, G1008, xenc228, G295, G306, G309, 
G334, xenc62, G359, G389, G1385, G1111, xenc11, G1165, G1267, G1886, 
G259, G262, G274, G296, xenc167, xenc45, G307, xenc202, G310, xenc97, 
G335, G360, G1242, xenc181, G390, G1828, G1868, G1869, xenc207, G1373, 
G1798, xenc37, xenc41, G1825, G265, G314, G336, xenc87, G407, G1293, 
G1294, G1892, xenc213, G1777, G1889, G410, xenc139, G1377, G1804, xenc188, 
G1237, G1829, G1295, G1670, G1678, G1729, G1737, G1761, G1769, xenc47, 
G340, G343, xenc156, G1781, G1238, xenc57, G1325, G1893, G1340, G1352, 
G1673, G1681, G1801, G1897, G1905, G391, G1299, xenc52, G1676, G1684, 
xenc134, G1081, G1733, xenc252, G1093, G1741, xenc26, G1765, G1773, G1239, 
xenc71, G1326, G1894, G1902, G392, G1360, xenc68, G1003, G1677, G1013, 
G1685, G1082, G1094, G1122, G1134, xenc10, G1187, G1805, G1327, G1901, 
xenc80, G1348, xenc19, G1909, G1758, G1766, xenc16, G377, G1243, G393, 
G1004, G1014, G1083, G1095, G1188, xenc98, G1900, xenc118, G1344, G1908, 
G1356, G1142, xenc216, G378, G399, G1331, G1005, G1015, G1764, G1126, 
G1130, G1772, G1138, xenc241, xenc112, G1189, G1343, xenc126, G1355, G324, 
G1099, xenc159, G379, G400, G449, G1087, G1088, G1125, xenc170, G1137, 
xenc247, G1345, xenc125, G1357, G1397, xenc35, G277, G1019, xenc6, G280, 
G1009, G325, xenc171, G364, G1193, xenc86, G401, xenc233, G1089, xenc39, 
G1127, xenc245, G1139, xenc163, G278, G281, xenc174, G326, G365, xenc76, 
G413, G1361, G1401, G445, G1349, G1350, G1389, G1493, G1501, xenc179, 
G1689, G279, G282, xenc107, G346, G1143, G366, G414, xenc135, G453, 
G1131, G1132, G1351, G1365, G1405, G285, xenc108, G347, xenc218, G367, 
G415, G1393, xenc104, G556, G1505, xenc120, G559, G1497, G1693, G1133, 
xenc90, G1477, G1485, xenc209, G1809, G348, G1369, G1409, G557, xenc49, 
G560, xenc150, G1362, G1378, G1429, G1437, G1686, G1774, xenc114, G1910, 
G1918, xenc32, xenc140, G544, G1489, G547, G1481, G558, xenc1, G561, 
G1813, G1370, G1368, xenc148, G417, G1384, G424, xenc238, G508, G1441, 
G511, G1433, G545, xenc21, G548, G564, G1692, G1024, G1780, G1148, 
G1916, xenc79, G1924, xenc146, G416, xenc196, G1376, G421, G423, G509, 
G512, xenc183, G546, xenc173, G549, G719, G722, G1023, G1147, xenc82, 
G418, xenc74, G420, G425, xenc65, G510, xenc116, G513, xenc110, G552, 
G1025, G1149, G419, xenc199, G422, xenc119, G441, G516, G725, G728, 
G1029, G1153, G433, G437, G663, G666, G731, G746, G756, G770, 
G1461, G1469, xenc38, G1413, G1421, G1445, G1453, G532, G1473, G535, 
G1465, xenc210, G495, G1425, G498, G1417, xenc182, G520, G1457, G523, 
G1449, G533, G536, xenc28, G496, G499, G521, xenc2, G524, xenc249, 
G534, xenc4, G537, G497, xenc103, G500, G522, G525, G540, G503, 
G528, G669, G672, xenc105, G569, G588, G618, xenc78, G639, G867, 
G588a, G588b, G639a, G639b, xenc93, G675, G688, G696, G710, xenc131, 
G73, G572, G573, G621, G622, xenc208, G776, G780, G784, G788, 
xenc24, G812, G832, G836, G1509, G1517, G1525, G1533, G1581, G1621, 
G1629, xenc73, G792, G796, G800, G804, G808, G816, G820, G824, 
G828, G871, G873, G875, G877, G879, G881, xenc158, G883, xenc194, 
G885, G1541, G1549, G1557, G1565, G1573, G1589, G1597, G1605, G1613, 
xenc193, G1, G1513, xenc31, G4, G1521, xenc164, G7, G1529, xenc235, 
G10, G1537, G28, G1585, xenc217, G43, G1625, xenc83, G46, G1633, 
xenc75, xenc133, G886, xenc160, G2, xenc129, G5, G8, G11, xenc48, 
G13, G1545, xenc219, xenc7, G16, G1553, G19, G1561, G22, G1569, 
G25, G1577, G29, G31, G1593, G34, G1601, G37, G1609, G40, 
G1617, G44, xenc89, G47, xenc72, xenc227, xenc55, G857, xenc46, xenc99, 
G860, G863, G865, xenc220, xenc166, xenc70, xenc153, xenc127, G14, xenc168, 
G17, xenc186, G20, G23, G26, G32, G35, xenc243, G38, G41, 
xenc88, xenc40, xenc198, G1913, G1921, xenc43, xenc232, xenc106, xenc221, xenc8, 
xenc204, xenc132, xenc63, xenc251, xenc214, G887, G462, xenc211, G74, G1637, 
G1917, xenc187, xenc225, G1647, G1925, xenc178, xenc58, G1020, G1144, G1386, 
G1394, G1402, G1638, G1648, G1806, xenc137, G1639, G1649, xenc157, G287, 
xenc56, G350, xenc192, G427, G429, xenc201, G431, G1028, G1152, G1392, 
G1400, G1408, G1812, xenc142, G1216, G286, G349, G426, xenc149, G428, 
G430, xenc51, G67, G1643, G70, G1653, G1215, G49, G53, G59, 
G61, G65, xenc234, G68, G71, xenc84, xenc226, G1217, xenc77, xenc34, 
xenc54, xenc180, xenc240, xenc253, xenc85, xenc189, xenc151, G375, G1221, G376, 
G55, xenc117;

not g0(G149, G101);
not g1(G153, G104);
not g2(G156, G107);
not g3(G160, G110);
not g4(G165, G113);
not g5(G168, G116);
not g6(G171, G119);
not g7(G175, G122);
not g8(G179, G125);
not g9(G184, G128);
not g10(G188, G131);
not g11(G191, G134);
not g12(G194, G137);
not g13(G198, G140);
not g14(G202, G143);
not g15(G206, G146);
nand g16(G231, G224, G898);
nand g17(G233, G227, G900);
not g18(G241, G237);
not g19(G244, G237);
assign G245 = G234;
assign G248 = G234;
not g22(G517, G469);
not g23(G529, G472);
not g24(G541, G475);
not g25(G553, G478);
not g26(G859, G953);
not g27(G862, G953);
not g28(G907, G898);
not g29(G909, G900);
assign G911 = G902;
not g31(G918, G902);
assign G919 = G902;
not g33(G922, G902);
assign G926 = G952;
not g35(G930, G952);
not g36(G932, G952);
assign G934 = G953;
not g38(G938, G953);
assign G943 = G953;
assign G947 = G953;
not g41(G949, G953);
assign G1506 = G101;
assign G1514 = G104;
assign G1522 = G107;
assign G1530 = G110;
assign G1538 = G113;
assign G1546 = G116;
assign G1554 = G119;
assign G1562 = G122;
assign G1570 = G125;
assign G1578 = G128;
assign G1586 = G131;
assign G1594 = G134;
assign G1602 = G137;
assign G1610 = G140;
assign G1618 = G143;
assign G1626 = G146;
not g58(G1512, G1506);
not g59(G1520, G1514);
not g60(G1528, G1522);
not g61(G1536, G1530);
not g62(G1544, G1538);
not g63(G1552, xenc200);
not g64(G1560, xenc231);
not g65(G1568, xenc33);
not g66(G1576, xenc14);
not g67(G1584, G1578);
not g68(G1592, xenc5);
not g69(G1600, G1594);
not g70(G1608, xenc9);
not g71(G1616, G1610);
not g72(G1624, xenc122);
not g73(G1632, G1626);
nand g74(G50, G930, xenc95);
nand g75(G52, G930, xenc95);
nand g76(G56, G930, xenc95);
nand g77(G58, G930, xenc95);
nand g78(G62, G930, xenc95);
nand g79(G64, G930, xenc95);
assign G251 = xenc169;
assign G254 = xenc100;
assign G288 = xenc124;
assign G291 = G168;
assign G299 = G184;
assign G302 = G202;
and g86(G318, G224, xenc0);
assign G321 = G179;
assign G327 = G188;
assign G330 = G191;
and g90(G352, G227, xenc0);
assign G355 = xenc244;
and g92(G369, G210, G241, xenc0);
assign G382 = xenc145;
assign G385 = xenc244;
nand g95(G853, xenc254, G907);
nand g96(G856, xenc254, G909);
nand g97(G893, xenc176, G237);
nand g98(G954, xenc176, xenc130);
nand g99(G955, G244, xenc130);
assign G1050 = xenc246;
assign G1053 = G175;
assign G1176 = G179;
assign G1179 = xenc244;
assign G1197 = xenc169;
assign G1207 = xenc169;
assign G1222 = xenc100;
assign G1244 = G188;
assign G1278 = G156;
and g109(G1290, G217, G245, xenc0);
assign G1300 = G191;
assign G1312 = xenc246;
assign G1332 = G194;
and g113(G1335, G221, G245, xenc0);
assign G1442 = G517;
assign G1450 = G517;
assign G1458 = G529;
assign G1466 = G529;
assign G1474 = G541;
assign G1482 = G541;
assign G1490 = xenc15;
assign G1498 = xenc15;
and g122(G1634, G231, G934);
and g123(G1644, G233, G934);
assign G1657 = G156;
assign G1665 = G156;
assign G1697 = xenc61;
assign G1705 = xenc61;
assign G1713 = xenc145;
assign G1721 = xenc145;
assign G1745 = G194;
assign G1753 = G194;
assign G1785 = xenc246;
assign G1793 = xenc246;
assign G1814 = xenc124;
assign G1817 = G175;
and g136(G1830, G214, G241, xenc0);
assign G1833 = G202;
assign G1841 = G179;
assign G1849 = G179;
assign G1854 = G168;
assign G1857 = G175;
assign G1870 = G184;
assign G1873 = G202;
assign G1878 = xenc61;
assign G1881 = G184;
not g146(G1642, G1634);
not g147(G1652, G1644);
not g148(G1056, G1050);
not g149(G1057, G1053);
not g150(G1182, G1176);
not g151(G1183, xenc60);
not g152(G1211, G1207);
not g153(G1298, xenc91);
not g154(G1320, G1312);
not g155(G1338, xenc111);
not g156(G1339, G1335);
and g157(G457, G210, xenc141);
and g158(G459, G217, xenc172);
nand g159(G482, G214, xenc141);
nand g160(G487, G221, xenc172);
nand g161(G492, G210, xenc141);
nand g162(G505, G217, xenc172);
not g163(G1456, G1450);
not g164(G1448, G1442);
not g165(G1472, xenc224);
not g166(G1464, G1458);
not g167(G1488, G1482);
not g168(G1480, xenc203);
not g169(G1504, G1498);
not g170(G1496, G1490);
nand g171(G956, G907, G919, xenc254, xenc184);
nand g172(G967, G909, G919, xenc254, xenc184);
nand g173(G978, G926, xenc212, xenc184);
and g174(G979, G926, xenc212, xenc184);
assign G980 = G251;
not g176(G1661, G1657);
assign G990 = G251;
not g178(G1669, G1665);
assign G1030 = G288;
not g180(G1701, xenc144);
assign G1040 = G288;
not g182(G1709, xenc152);
assign G1058 = G299;
not g184(G1717, G1713);
assign G1068 = G299;
not g186(G1725, G1721);
assign G1078 = xenc197;
assign G1090 = xenc197;
assign G1100 = G327;
not g190(G1749, G1745);
assign G1112 = G327;
not g192(G1757, xenc59);
assign G1154 = G352;
not g194(G1789, xenc223);
assign G1166 = G352;
not g196(G1797, G1793);
assign G1194 = xenc67;
not g198(G1201, G1197);
assign G1204 = xenc67;
not g200(G1820, xenc36);
not g201(G1821, G1817);
not g202(G1230, xenc229);
not g203(G1836, xenc94);
not g204(G1837, G1833);
not g205(G1252, G1244);
assign G1256 = G382;
not g207(G1845, G1841);
assign G1268 = G382;
not g209(G1853, G1849);
not g210(G1860, xenc239);
not g211(G1861, G1857);
not g212(G1286, G1278);
not g213(G1876, G1870);
not g214(G1877, G1873);
not g215(G1308, G1300);
not g216(G1884, xenc44);
not g217(G1885, G1881);
assign G1654 = xenc12;
assign G1662 = xenc12;
assign G1694 = G291;
assign G1702 = G291;
assign G1710 = xenc29;
assign G1718 = xenc29;
assign G1726 = G321;
assign G1734 = G321;
assign G1742 = G330;
assign G1750 = G330;
assign G1782 = G355;
assign G1790 = G355;
assign G1838 = G385;
assign G1846 = G385;
nand g232(G297, G1053, xenc250);
nand g233(G298, G1050, xenc3);
nand g234(G361, xenc60, G1182);
nand g235(G362, G1176, xenc206);
nand g236(G404, G1335, xenc162);
nand g237(G405, xenc111, G1339);
nand g238(G1225, G1817, G1820);
nand g239(G1226, xenc36, G1821);
nand g240(G1247, G1833, G1836);
nand g241(G1248, xenc94, xenc165);
nand g242(G1281, G1857, G1860);
nand g243(G1282, xenc239, G1861);
nand g244(G1303, G1873, xenc190);
nand g245(G1304, G1870, G1877);
nand g246(G1315, G1881, G1884);
nand g247(G1316, xenc44, xenc154);
not g248(G998, xenc155);
not g249(G988, G980);
nand g250(G268, G297, G298);
not g251(G1038, G1030);
not g252(G1048, G1040);
not g253(G1076, G1068);
not g254(G1066, G1058);
not g255(G1098, G1090);
not g256(G1120, xenc195);
not g257(G1174, G1166);
nand g258(G363, G361, G362);
not g259(G1210, G1204);
nand g260(G373, G1204, G1211);
not g261(G1276, G1268);
nand g262(G406, xenc161, G405);
not g263(G565, G482);
assign G566 = G482;
not g265(G614, G487);
assign G615 = G487;
nand g267(G958, G956, G978);
nand g268(G969, G967, G978);
not g269(G1660, xenc147);
nand g270(G984, xenc147, xenc255);
not g271(G1668, G1662);
nand g272(G994, G1662, G1669);
not g273(G1700, G1694);
nand g274(G1034, G1694, xenc191);
not g275(G1708, G1702);
nand g276(G1044, G1702, xenc138);
not g277(G1716, xenc27);
nand g278(G1062, xenc27, G1717);
not g279(G1724, G1718);
nand g280(G1072, G1718, G1725);
not g281(G1732, G1726);
not g282(G1086, xenc121);
not g283(G1740, G1734);
not g284(G1748, xenc53);
nand g285(G1104, xenc53, xenc177);
not g286(G1108, xenc25);
not g287(G1756, G1750);
nand g288(G1116, G1750, xenc96);
not g289(G1788, G1782);
nand g290(G1158, G1782, G1789);
not g291(G1162, G1154);
not g292(G1796, G1790);
nand g293(G1170, G1790, G1797);
not g294(G1200, G1194);
nand g295(G1203, G1194, G1201);
nand g296(G1227, G1225, G1226);
nand g297(G1249, G1247, G1248);
not g298(G1844, G1838);
nand g299(G1260, G1838, G1845);
not g300(G1264, G1256);
not g301(G1852, G1846);
nand g302(G1272, G1846, G1853);
nand g303(G1283, G1281, xenc113);
nand g304(G1305, xenc20, xenc69);
nand g305(G1317, G1315, G1316);
assign G1410 = G492;
assign G1418 = G492;
assign G1426 = xenc17;
assign G1434 = xenc17;
not g310(G269, xenc222);
nand g311(G372, G1207, xenc185);
nand g312(G983, G1657, xenc205);
nand g313(G993, G1665, G1668);
nand g314(G1033, xenc144, G1700);
nand g315(G1043, xenc152, G1708);
nand g316(G1061, G1713, G1716);
nand g317(G1071, G1721, G1724);
nand g318(G1103, G1745, G1748);
nand g319(G1115, xenc59, G1756);
nand g320(G1157, xenc223, xenc237);
nand g321(G1169, G1793, G1796);
not g322(G1184, xenc101);
nand g323(G1202, G1197, G1200);
nand g324(G1259, G1841, G1844);
nand g325(G1271, G1849, G1852);
not g326(G1322, G406);
nand g327(G374, G372, xenc248);
nand g328(G396, xenc230, xenc102);
not g329(G1321, xenc230);
not g330(G1424, G1418);
not g331(G1416, G1410);
not g332(G1440, G1434);
not g333(G1432, G1426);
nand g334(G985, G983, xenc242);
nand g335(G995, G993, G994);
nand g336(G1035, G1033, G1034);
nand g337(G1045, G1043, G1044);
nand g338(G1063, G1061, xenc175);
nand g339(G1073, G1071, G1072);
nand g340(G1105, G1103, xenc23);
nand g341(G1117, xenc50, G1116);
nand g342(G1159, G1157, G1158);
nand g343(G1171, G1169, G1170);
nand g344(G1212, G1202, G1203);
not g345(G1231, G1227);
nand g346(G1232, G1227, G1230);
not g347(G1253, G1249);
nand g348(G1254, G1249, xenc236);
nand g349(G1261, G1259, G1260);
nand g350(G1273, xenc64, xenc109);
not g351(G1287, G1283);
nand g352(G1288, G1283, G1286);
not g353(G1309, G1305);
nand g354(G1310, G1305, G1308);
not g355(G1192, G1184);
nand g356(G397, G1312, G1321);
not g357(G1330, G1322);
assign G1000 = G269;
assign G1010 = G269;
nand g360(G1233, xenc229, G1231);
nand g361(G1255, G1244, G1253);
nand g362(G1289, G1278, xenc18);
nand g363(G1311, G1300, xenc136);
not g364(G1381, G374);
nand g365(G257, G995, G998);
not g366(G999, G995);
nand g367(G260, G985, G988);
not g368(G989, G985);
nand g369(G272, G1035, G1038);
not g370(G1039, G1035);
nand g371(G294, G1045, G1048);
not g372(G1049, G1045);
nand g373(G305, G1073, G1076);
not g374(G1077, G1073);
nand g375(G308, G1063, xenc128);
not g376(G1067, G1063);
nand g377(G333, xenc22, xenc42);
not g378(G1121, xenc22);
nand g379(G358, G1171, G1174);
not g380(G1175, G1171);
not g381(G1220, xenc143);
nand g382(G388, xenc66, xenc123);
not g383(G1277, xenc66);
nand g384(G398, G396, G397);
not g385(G1109, xenc215);
nand g386(G1110, xenc215, G1108);
not g387(G1163, xenc30);
nand g388(G1164, xenc30, G1162);
nand g389(G1234, G1232, G1233);
not g390(G1265, G1261);
nand g391(G1266, G1261, G1264);
nand g392(G1822, G1254, G1255);
nand g393(G1862, G1310, G1311);
nand g394(G1865, xenc115, G1289);
nand g395(G258, xenc155, xenc92);
nand g396(G261, G980, xenc81);
nand g397(G273, G1030, G1039);
not g398(G1018, xenc13);
not g399(G1008, G1000);
nand g400(G295, G1040, xenc228);
nand g401(G306, G1068, G1077);
nand g402(G309, G1058, G1067);
nand g403(G334, xenc195, G1121);
nand g404(G359, G1166, xenc62);
nand g405(G389, G1268, G1277);
not g406(G1385, G1381);
nand g407(G1111, xenc25, G1109);
nand g408(G1165, G1154, xenc11);
nand g409(G1267, G1256, G1265);
not g410(G1886, G398);
nand g411(G259, G257, G258);
nand g412(G262, G260, G261);
nand g413(G274, G272, G273);
nand g414(G296, G294, G295);
nand g415(G307, xenc167, xenc45);
nand g416(G310, xenc202, G309);
nand g417(G335, G333, xenc97);
nand g418(G360, G358, G359);
not g419(G1242, G1234);
nand g420(G390, xenc181, G389);
not g421(G1828, G1822);
not g422(G1868, G1862);
not g423(G1869, G1865);
nand g424(G1373, G1164, xenc207);
nand g425(G1798, G1110, G1111);
nand g426(G1825, xenc37, xenc41);
not g427(G265, G259);
not g428(G314, G307);
not g429(G336, G335);
not g430(G407, xenc87);
nand g431(G1293, G1865, G1868);
nand g432(G1294, G1862, G1869);
not g433(G1892, G1886);
not g434(G1777, xenc213);
not g435(G1889, G390);
assign G410 = G310;
not g437(G1377, xenc139);
not g438(G1804, G1798);
nand g439(G1237, G1825, xenc188);
not g440(G1829, G1825);
nand g441(G1295, G1293, G1294);
assign G1670 = G274;
assign G1678 = G274;
assign G1729 = G310;
assign G1737 = G310;
assign G1761 = G262;
assign G1769 = G262;
assign G340 = xenc47;
assign G343 = G314;
not g450(G1781, xenc156);
nand g451(G1238, G1822, G1829);
nand g452(G1325, xenc57, G1892);
not g453(G1893, xenc57);
assign G1340 = G407;
assign G1352 = G407;
assign G1673 = G265;
assign G1681 = G265;
assign G1801 = G314;
assign G1897 = xenc47;
assign G1905 = xenc47;
nand g461(G391, G1295, G1298);
not g462(G1299, G1295);
not g463(G1676, xenc52);
not g464(G1684, G1678);
nand g465(G1081, G1729, xenc134);
not g466(G1733, G1729);
nand g467(G1093, G1737, xenc252);
not g468(G1741, G1737);
not g469(G1765, xenc26);
not g470(G1773, G1769);
nand g471(G1239, G1237, G1238);
nand g472(G1326, G1886, xenc71);
assign G1894 = G410;
assign G1902 = G410;
nand g475(G392, xenc91, G1299);
not g476(G1360, G1352);
nand g477(G1003, G1673, xenc68);
not g478(G1677, G1673);
nand g479(G1013, G1681, G1684);
not g480(G1685, G1681);
nand g481(G1082, G1726, G1733);
nand g482(G1094, G1734, G1741);
assign G1122 = G340;
assign G1134 = G340;
nand g485(G1187, xenc10, G1804);
not g486(G1805, xenc10);
nand g487(G1327, G1325, G1326);
not g488(G1901, G1897);
not g489(G1348, xenc80);
not g490(G1909, xenc19);
assign G1758 = G343;
assign G1766 = G343;
nand g493(G377, G1239, xenc16);
not g494(G1243, G1239);
nand g495(G393, G391, G392);
nand g496(G1004, xenc52, G1677);
nand g497(G1014, G1678, G1685);
nand g498(G1083, G1081, G1082);
nand g499(G1095, G1093, G1094);
nand g500(G1188, G1798, G1805);
not g501(G1900, xenc98);
nand g502(G1344, xenc98, xenc118);
not g503(G1908, G1902);
nand g504(G1356, G1902, G1909);
not g505(G1142, G1134);
nand g506(G378, G1234, xenc216);
nand g507(G399, G1327, G1330);
not g508(G1331, G1327);
nand g509(G1005, G1003, G1004);
nand g510(G1015, G1013, G1014);
not g511(G1764, G1758);
nand g512(G1126, G1758, G1765);
not g513(G1130, G1122);
not g514(G1772, G1766);
nand g515(G1138, G1766, G1773);
nand g516(G1189, xenc241, xenc112);
nand g517(G1343, G1897, G1900);
nand g518(G1355, xenc19, xenc126);
nand g519(G324, G1095, G1098);
not g520(G1099, G1095);
nand g521(G379, xenc159, G378);
nand g522(G400, G1322, G1331);
nand g523(G449, G393, G918);
not g524(G1087, G1083);
nand g525(G1088, G1083, G1086);
nand g526(G1125, xenc26, G1764);
nand g527(G1137, G1769, xenc170);
nand g528(G1345, xenc247, G1344);
nand g529(G1357, xenc125, G1356);
assign G1397 = G393;
nand g531(G277, xenc35, G1018);
not g532(G1019, xenc35);
nand g533(G280, G1005, xenc6);
not g534(G1009, G1005);
nand g535(G325, G1090, G1099);
nand g536(G364, G1189, xenc171);
not g537(G1193, G1189);
nand g538(G401, G399, xenc86);
nand g539(G1089, xenc121, xenc233);
nand g540(G1127, G1125, xenc39);
nand g541(G1139, xenc245, G1138);
nand g542(G278, xenc13, xenc163);
nand g543(G281, G1000, G1009);
nand g544(G326, G324, xenc174);
nand g545(G365, G1184, G1193);
nand g546(G413, G1357, xenc76);
not g547(G1361, G1357);
not g548(G1401, G1397);
nand g549(G445, G379, G918);
not g550(G1349, G1345);
nand g551(G1350, G1345, G1348);
assign G1389 = G379;
assign G1493 = G449;
assign G1501 = G449;
nand g555(G1689, xenc179, G1089);
nand g556(G279, G277, G278);
nand g557(G282, G280, G281);
nand g558(G346, xenc107, G1142);
not g559(G1143, xenc107);
nand g560(G366, G364, G365);
nand g561(G414, G1352, G1361);
nand g562(G453, xenc135, G918);
not g563(G1131, G1127);
nand g564(G1132, G1127, G1130);
nand g565(G1351, xenc80, G1349);
not g566(G1365, G326);
assign G1405 = xenc135;
not g568(G285, G279);
nand g569(G347, G1134, xenc108);
not g570(G367, xenc218);
nand g571(G415, G413, G414);
not g572(G1393, G1389);
nand g573(G556, G1501, xenc104);
not g574(G1505, G1501);
nand g575(G559, G1493, xenc120);
not g576(G1497, G1493);
not g577(G1693, G1689);
nand g578(G1133, G1122, G1131);
assign G1477 = xenc90;
assign G1485 = xenc90;
nand g581(G1809, G1350, xenc209);
nand g582(G348, G346, G347);
not g583(G1369, G1365);
not g584(G1409, G1405);
nand g585(G557, G1498, G1505);
nand g586(G560, G1490, xenc49);
assign G1362 = xenc150;
not g588(G1378, G415);
assign G1429 = G453;
assign G1437 = G453;
assign G1686 = xenc150;
nand g592(G1774, G1132, G1133);
and g593(G1910, G285, xenc114);
and g594(G1918, G856, G367);
nand g595(G544, xenc32, xenc140);
not g596(G1489, xenc32);
nand g597(G547, G1477, G1480);
not g598(G1481, G1477);
nand g599(G558, G556, G557);
nand g600(G561, G559, xenc1);
not g601(G1813, G1809);
not g602(G1370, G348);
not g603(G1368, G1362);
nand g604(G417, G1362, xenc148);
not g605(G1384, G1378);
nand g606(G424, G1378, G1385);
nand g607(G508, xenc238, G1440);
not g608(G1441, xenc238);
nand g609(G511, G1429, G1432);
not g610(G1433, G1429);
nand g611(G545, G1482, G1489);
nand g612(G548, xenc203, xenc21);
not g613(G564, G558);
not g614(G1692, G1686);
nand g615(G1024, G1686, G1693);
not g616(G1780, G1774);
nand g617(G1148, G1774, G1781);
not g618(G1916, G1910);
not g619(G1924, xenc79);
nand g620(G416, G1365, xenc146);
not g621(G1376, xenc196);
nand g622(G421, xenc196, G1377);
nand g623(G423, G1381, G1384);
nand g624(G509, G1434, G1441);
nand g625(G512, G1426, G1433);
nand g626(G546, G544, xenc183);
nand g627(G549, G547, xenc173);
not g628(G719, G561);
assign G722 = G561;
nand g630(G1023, G1689, G1692);
nand g631(G1147, xenc156, G1780);
nand g632(G418, G416, xenc82);
nand g633(G420, xenc139, xenc74);
nand g634(G425, G423, G424);
nand g635(G510, xenc65, G509);
nand g636(G513, xenc116, G512);
not g637(G552, xenc110);
nand g638(G1025, G1023, G1024);
nand g639(G1149, G1147, G1148);
not g640(G419, G418);
nand g641(G422, xenc199, G421);
nand g642(G441, xenc119, G918);
not g643(G516, G510);
not g644(G725, G549);
assign G728 = G549;
not g646(G1029, G1025);
not g647(G1153, G1149);
nand g648(G433, G419, G918);
nand g649(G437, G422, G918);
not g650(G663, G513);
assign G666 = G513;
and g652(G731, G719, G725);
and g653(G746, G722, G725);
and g654(G756, G719, G728);
and g655(G770, G722, G728);
assign G1461 = G441;
assign G1469 = G441;
assign G1413 = xenc38;
assign G1421 = xenc38;
assign G1445 = G437;
assign G1453 = G437;
nand g662(G532, G1469, G1472);
not g663(G1473, G1469);
nand g664(G535, G1461, G1464);
not g665(G1465, G1461);
nand g666(G495, G1421, xenc210);
not g667(G1425, G1421);
nand g668(G498, G1413, G1416);
not g669(G1417, G1413);
nand g670(G520, G1453, xenc182);
not g671(G1457, G1453);
nand g672(G523, G1445, G1448);
not g673(G1449, G1445);
nand g674(G533, xenc224, G1473);
nand g675(G536, G1458, G1465);
nand g676(G496, G1418, xenc28);
nand g677(G499, G1410, G1417);
nand g678(G521, G1450, G1457);
nand g679(G524, G1442, xenc2);
nand g680(G534, xenc249, G533);
nand g681(G537, xenc4, G536);
nand g682(G497, G495, G496);
nand g683(G500, xenc103, G499);
nand g684(G522, G520, G521);
nand g685(G525, G523, G524);
not g686(G540, G534);
not g687(G503, G497);
not g688(G528, G522);
not g689(G669, G537);
assign G672 = G537;
not g691(G569, xenc105);
and g692(G588, G566, xenc105);
not g693(G618, G525);
and g694(G639, xenc78, G525);
nand g695(G867, G516, G564, G552, G540, G482, G528, G503, G487);
assign G588a = G588;
assign G588b = G588;
assign G639a = G639;
assign G639b = G639;
and g700(G675, xenc93, G669);
and g701(G688, G666, G669);
and g702(G696, xenc93, G672);
and g703(G710, G666, G672);
and g704(G73, xenc212, G867, xenc131, xenc131);
and g705(G572, G565, G569);
and g706(G573, G566, G569);
and g707(G621, G614, G618);
and g708(G622, xenc78, G618);
nand g709(G776, G588a, G639a, G696, xenc208, G958);
nand g710(G780, G588a, G639a, G675, G756, G958);
nand g711(G784, G588a, G639a, G675, G746, G958);
nand g712(G788, G588a, G639a, G688, xenc208, G958);
nand g713(G812, G588b, G639a, xenc24, G746, G969);
nand g714(G832, G588b, G639b, G696, G770, G969);
nand g715(G836, G588b, G639b, xenc24, G756, G969);
and g716(G1509, G588a, G639a, G696, xenc208, G958);
and g717(G1517, G588a, G639a, G675, G756, G958);
and g718(G1525, G588a, G639a, G675, G746, G958);
and g719(G1533, G588a, G639a, G688, xenc208, G958);
and g720(G1581, G588b, G639a, xenc24, G746, G969);
and g721(G1621, G588b, G639b, G696, G770, G969);
and g722(G1629, G588b, G639b, xenc24, G756, G969);
nand g723(G792, G588a, xenc73, G696, G756, G958);
nand g724(G796, G588b, xenc73, G696, G746, G958);
nand g725(G800, G588b, xenc73, xenc24, xenc208, G958);
nand g726(G804, G588b, xenc73, G675, G770, G958);
nand g727(G808, G588b, xenc73, G688, G756, G969);
nand g728(G816, G573, G639b, G696, G756, G969);
nand g729(G820, G573, G639b, G696, G746, G969);
nand g730(G824, G573, G639b, xenc24, xenc208, G969);
nand g731(G828, G573, G639b, G688, G756, G969);
nand g732(G871, G588b, xenc73, G675, xenc208, G979);
nand g733(G873, G573, G639b, G675, xenc208, G979);
nand g734(G875, G573, xenc73, G696, xenc208, G979);
nand g735(G877, G573, xenc73, G675, G756, G979);
nand g736(G879, G573, xenc73, G675, G746, G979);
nand g737(G881, G573, xenc73, G688, xenc208, G979);
nand g738(G883, G573, xenc158, G675, xenc208, G979);
nand g739(G885, xenc194, xenc73, G675, xenc208, G979);
and g740(G1541, G588a, xenc73, G696, G756, G958);
and g741(G1549, G588b, xenc73, G696, G746, G958);
and g742(G1557, G588b, xenc73, xenc24, xenc208, G958);
and g743(G1565, G588b, xenc73, G675, G770, G958);
and g744(G1573, G588b, xenc73, G688, G756, G969);
and g745(G1589, G573, G639b, G696, G756, G969);
and g746(G1597, G573, G639b, G696, G746, G969);
and g747(G1605, G573, G639b, xenc24, xenc208, G969);
and g748(G1613, G573, G639b, G688, G756, G969);
nand g749(G1, G1509, xenc193);
not g750(G1513, G1509);
nand g751(G4, G1517, xenc31);
not g752(G1521, G1517);
nand g753(G7, xenc164, G1528);
not g754(G1529, xenc164);
nand g755(G10, xenc235, G1536);
not g756(G1537, xenc235);
nand g757(G28, G1581, G1584);
not g758(G1585, G1581);
nand g759(G43, xenc217, G1624);
not g760(G1625, xenc217);
nand g761(G46, xenc83, G1632);
not g762(G1633, xenc83);
and g763(G886, G871, xenc75, G875, G877, G879, G881, xenc133, G885);
nand g764(G2, G1506, xenc160);
nand g765(G5, G1514, xenc129);
nand g766(G8, G1522, G1529);
nand g767(G11, G1530, G1537);
nand g768(G13, G1541, xenc48);
not g769(G1545, G1541);
nand g770(G16, xenc219, xenc7);
not g771(G1553, xenc219);
nand g772(G19, G1557, G1560);
not g773(G1561, G1557);
nand g774(G22, G1565, G1568);
not g775(G1569, G1565);
nand g776(G25, G1573, G1576);
not g777(G1577, G1573);
nand g778(G29, G1578, G1585);
nand g779(G31, G1589, G1592);
not g780(G1593, G1589);
nand g781(G34, G1597, G1600);
not g782(G1601, G1597);
nand g783(G37, G1605, G1608);
not g784(G1609, G1605);
nand g785(G40, G1613, G1616);
not g786(G1617, G1613);
nand g787(G44, xenc122, G1625);
nand g788(G47, G1626, xenc89);
nand g789(G857, G776, xenc72, G784, xenc227, G792, xenc55, G800, G804);
nand g790(G860, G808, G812, xenc46, G820, xenc99, G828, G832, G836);
and g791(G863, G776, xenc72, G784, xenc227, G792, xenc55, G800, G804);
and g792(G865, G808, G812, xenc46, G820, xenc99, G828, G832, G836);
nand g793(xenc166, G1, xenc220);
nand g794(xenc70, G4, G5);
nand g795(G9, G7, xenc153);
nand g796(xenc127, G10, G11);
nand g797(G14, G1538, G1545);
nand g798(G17, xenc200, xenc168);
nand g799(G20, xenc231, xenc186);
nand g800(G23, xenc33, G1569);
nand g801(G26, xenc14, G1577);
nand g802(G30, G28, G29);
nand g803(G32, xenc5, G1593);
nand g804(G35, G1594, G1601);
nand g805(G38, xenc9, xenc243);
nand g806(G41, G1610, G1617);
nand g807(xenc40, G43, xenc88);
nand g808(xenc198, G46, G47);
and g809(G1913, G857, G859);
and g810(G1921, G860, G862);
nand g811(G15, G13, G14);
nand g812(G18, xenc43, G17);
nand g813(xenc232, G19, G20);
nand g814(G24, G22, xenc106);
nand g815(xenc221, G25, G26);
nand g816(xenc8, G31, G32);
nand g817(G36, G34, G35);
nand g818(xenc63, xenc204, xenc132);
nand g819(G42, xenc251, xenc214);
and g820(G887, G863, G865, G886);
nand g821(G462, G863, G865);
and g822(G74, xenc212, G867, G952, xenc211);
nand g823(G1637, G1913, G1916);
not g824(G1917, G1913);
nand g825(G1647, xenc187, xenc225);
not g826(G1925, xenc187);
nor g827(G75, xenc178, G74);
and g828(G1020, G457, G911, xenc58);
and g829(G1144, G469, G911, xenc58);
and g830(G1386, G475, G911, xenc58);
and g831(G1394, G478, G911, xenc58);
and g832(G1402, G459, G911, xenc58);
nand g833(G1638, G1910, G1917);
nand g834(G1648, xenc79, G1925);
and g835(G1806, G472, G911, xenc58);
nand g836(G1639, G1637, xenc137);
nand g837(G1649, G1647, G1648);
nand g838(G287, xenc157, G1029);
nand g839(G350, xenc56, G1153);
nand g840(G427, G1386, xenc192);
nand g841(G429, G1394, G1401);
nand g842(G431, xenc201, G1409);
not g843(G1028, xenc157);
not g844(G1152, xenc56);
not g845(G1392, G1386);
not g846(G1400, G1394);
not g847(G1408, xenc201);
not g848(G1812, G1806);
nand g849(G1216, G1806, xenc142);
nand g850(G286, G1025, G1028);
nand g851(G349, G1149, G1152);
nand g852(G426, G1389, G1392);
nand g853(G428, G1397, xenc149);
nand g854(G430, G1405, G1408);
nand g855(G67, xenc51, G1642);
not g856(G1643, xenc51);
nand g857(G70, G1649, G1652);
not g858(G1653, G1649);
nand g859(G1215, G1809, G1812);
nand g860(G49, G286, G287);
nand g861(G53, G349, G350);
nand g862(G59, G426, G427);
nand g863(G61, G428, G429);
nand g864(G65, G430, G431);
nand g865(G68, G1634, xenc234);
nand g866(G71, G1644, G1653);
nand g867(G1217, xenc84, xenc226);
and g868(xenc34, G49, xenc77);
and g869(xenc180, G52, xenc54);
and g870(G60, xenc240, xenc253);
and g871(G63, G61, G62);
and g872(G66, xenc85, xenc189);
nand g873(xenc151, G67, G68);
nand g874(G72, G70, G71);
nand g875(G375, G1217, G1220);
not g876(G1221, G1217);
nand g877(G376, xenc143, G1221);
nand g878(G55, G375, G376);
and g879(G57, xenc117, G56);
xnor g880(xenc0, G938, keyinput0);
xnor g881(xenc1, G560, keyinput1);
xnor g882(xenc2, G1449, keyinput2);
xor g883(xenc3, G1057, keyinput3);
xor g884(xenc4, G535, keyinput4);
xor g885(xenc5, G1586, keyinput5);
xnor g886(xenc6, G1008, keyinput6);
xnor g887(xenc7, G1552, keyinput7);
xnor g888(G33, xenc8, keyinput8);
xor g889(xenc9, G1602, keyinput9);
xnor g890(xenc10, G1801, keyinput10);
xor g891(xenc11, G1163, keyinput11);
xnor g892(xenc12, G254, keyinput12);
xnor g893(xenc13, G1010, keyinput13);
xor g894(xenc14, G1570, keyinput14);
xor g895(xenc15, G553, keyinput15);
xnor g896(xenc16, G1242, keyinput16);
xor g897(xenc17, G505, keyinput17);
xnor g898(xenc18, G1287, keyinput18);
xnor g899(xenc19, G1905, keyinput19);
xnor g900(xenc20, G1303, keyinput20);
xnor g901(xenc21, G1481, keyinput21);
xnor g902(xenc22, G1117, keyinput22);
xnor g903(xenc23, G1104, keyinput23);
xnor g904(xenc24, G710, keyinput24);
xnor g905(xenc25, G1100, keyinput25);
xnor g906(xenc26, G1761, keyinput26);
xor g907(xenc27, G1710, keyinput27);
xor g908(xenc28, G1425, keyinput28);
xor g909(xenc29, G302, keyinput29);
xor g910(xenc30, G1159, keyinput30);
xor g911(xenc31, G1520, keyinput31);
xnor g912(xenc32, G1485, keyinput32);
xor g913(xenc33, G1562, keyinput33);
xnor g914(G51, xenc34, keyinput34);
xor g915(xenc35, G1015, keyinput35);
xor g916(xenc36, G1814, keyinput36);
xnor g917(xenc37, G1266, keyinput37);
xnor g918(xenc38, G433, keyinput38);
xor g919(xenc39, G1126, keyinput39);
xor g920(G45, xenc40, keyinput40);
xnor g921(xenc41, G1267, keyinput41);
xnor g922(xenc42, G1120, keyinput42);
xor g923(xenc43, G16, keyinput43);
xnor g924(xenc44, G1878, keyinput44);
xnor g925(xenc45, G306, keyinput45);
xor g926(xenc46, G816, keyinput46);
xnor g927(xenc47, G336, keyinput47);
xor g928(xenc48, G1544, keyinput48);
xor g929(xenc49, G1497, keyinput49);
xnor g930(xenc50, G1115, keyinput50);
xnor g931(xenc51, G1639, keyinput51);
xor g932(xenc52, G1670, keyinput52);
xor g933(xenc53, G1742, keyinput53);
xnor g934(xenc54, G53, keyinput54);
xor g935(xenc55, G796, keyinput55);
xor g936(xenc56, G1144, keyinput56);
xor g937(xenc57, G1889, keyinput57);
xor g938(xenc58, G462, keyinput58);
xnor g939(xenc59, G1753, keyinput59);
xnor g940(xenc60, G1179, keyinput60);
xnor g941(xenc61, G171, keyinput61);
xnor g942(xenc62, G1175, keyinput62);
xnor g943(G39, xenc63, keyinput63);
xnor g944(xenc64, G1271, keyinput64);
xnor g945(xenc65, G508, keyinput65);
xnor g946(xenc66, G1273, keyinput66);
xor g947(xenc67, G369, keyinput67);
xor g948(xenc68, G1676, keyinput68);
xnor g949(xenc69, G1304, keyinput69);
xnor g950(G6, xenc70, keyinput70);
xnor g951(xenc71, G1893, keyinput71);
xnor g952(xenc72, G780, keyinput72);
xnor g953(xenc73, G622, keyinput73);
xnor g954(xenc74, G1376, keyinput74);
xnor g955(xenc75, G873, keyinput75);
xnor g956(xenc76, G1360, keyinput76);
xor g957(xenc77, G50, keyinput77);
xnor g958(xenc78, G615, keyinput78);
xnor g959(xenc79, G1918, keyinput79);
xnor g960(xenc80, G1340, keyinput80);
xnor g961(xenc81, G989, keyinput81);
xnor g962(xenc82, G417, keyinput82);
xor g963(xenc83, G1629, keyinput83);
xor g964(xenc84, G1215, keyinput84);
xnor g965(xenc85, G64, keyinput85);
xnor g966(xenc86, G400, keyinput86);
xnor g967(xenc87, G296, keyinput87);
xor g968(xenc88, G44, keyinput88);
xor g969(xenc89, G1633, keyinput89);
xor g970(xenc90, G445, keyinput90);
xnor g971(xenc91, G1290, keyinput91);
xnor g972(xenc92, G999, keyinput92);
xor g973(xenc93, G663, keyinput93);
xnor g974(xenc94, G1830, keyinput94);
xnor g975(xenc95, G947, keyinput95);
xor g976(xenc96, G1757, keyinput96);
xnor g977(xenc97, G334, keyinput97);
xor g978(xenc98, G1894, keyinput98);
xnor g979(xenc99, G824, keyinput99);
xnor g980(xenc100, G153, keyinput100);
xor g981(xenc101, G363, keyinput101);
xor g982(xenc102, G1320, keyinput102);
xnor g983(xenc103, G498, keyinput103);
xor g984(xenc104, G1504, keyinput104);
xor g985(xenc105, G500, keyinput105);
xnor g986(xenc106, G23, keyinput106);
xnor g987(xenc107, G1139, keyinput107);
xnor g988(xenc108, G1143, keyinput108);
xnor g989(xenc109, G1272, keyinput109);
xnor g990(xenc110, G546, keyinput110);
xnor g991(xenc111, G1332, keyinput111);
xor g992(xenc112, G1188, keyinput112);
xnor g993(xenc113, G1282, keyinput113);
xor g994(xenc114, G853, keyinput114);
xnor g995(xenc115, G1288, keyinput115);
xnor g996(xenc116, G511, keyinput116);
xor g997(xenc117, G55, keyinput117);
xor g998(xenc118, G1901, keyinput118);
xnor g999(xenc119, G425, keyinput119);
xor g1000(xenc120, G1496, keyinput120);
xnor g1001(xenc121, G1078, keyinput121);
xnor g1002(xenc122, G1618, keyinput122);
xor g1003(xenc123, G1276, keyinput123);
xor g1004(xenc124, G165, keyinput124);
xnor g1005(xenc125, G1355, keyinput125);
xor g1006(xenc126, G1908, keyinput126);
xnor g1007(G12, xenc127, keyinput127);
xor g1008(xenc128, G1066, keyinput128);
xnor g1009(xenc129, G1521, keyinput129);
xor g1010(xenc130, G922, keyinput130);
xor g1011(xenc131, G932, keyinput131);
xor g1012(xenc132, G38, keyinput132);
xnor g1013(xenc133, G883, keyinput133);
xnor g1014(xenc134, G1732, keyinput134);
xnor g1015(xenc135, G401, keyinput135);
xor g1016(xenc136, G1309, keyinput136);
xnor g1017(xenc137, G1638, keyinput137);
xnor g1018(xenc138, G1709, keyinput138);
xor g1019(xenc139, G1373, keyinput139);
xor g1020(xenc140, G1488, keyinput140);
xnor g1021(xenc141, G955, keyinput141);
xor g1022(xenc142, G1813, keyinput142);
xnor g1023(xenc143, G1212, keyinput143);
xnor g1024(xenc144, G1697, keyinput144);
xnor g1025(xenc145, G206, keyinput145);
xnor g1026(xenc146, G1368, keyinput146);
xor g1027(xenc147, G1654, keyinput147);
xor g1028(xenc148, G1369, keyinput148);
xor g1029(xenc149, G1400, keyinput149);
xor g1030(xenc150, G282, keyinput150);
xnor g1031(G69, xenc151, keyinput151);
xor g1032(xenc152, G1705, keyinput152);
xor g1033(xenc153, G8, keyinput153);
xor g1034(xenc154, G1885, keyinput154);
xnor g1035(xenc155, G990, keyinput155);
xor g1036(xenc156, G1777, keyinput156);
xnor g1037(xenc157, G1020, keyinput157);
xor g1038(xenc158, G621, keyinput158);
xnor g1039(xenc159, G377, keyinput159);
xnor g1040(xenc160, G1513, keyinput160);
xnor g1041(xenc161, G404, keyinput161);
xnor g1042(xenc162, G1338, keyinput162);
xor g1043(xenc163, G1019, keyinput163);
xnor g1044(xenc164, G1525, keyinput164);
xnor g1045(xenc165, G1837, keyinput165);
xnor g1046(G3, xenc166, keyinput166);
xor g1047(xenc167, G305, keyinput167);
xnor g1048(xenc168, G1553, keyinput168);
xnor g1049(xenc169, G149, keyinput169);
xnor g1050(xenc170, G1772, keyinput170);
xor g1051(xenc171, G1192, keyinput171);
xor g1052(xenc172, G954, keyinput172);
xor g1053(xenc173, G548, keyinput173);
xor g1054(xenc174, G325, keyinput174);
xor g1055(xenc175, G1062, keyinput175);
xor g1056(xenc176, G248, keyinput176);
xnor g1057(xenc177, G1749, keyinput177);
xnor g1058(xenc178, G73, keyinput178);
xnor g1059(xenc179, G1088, keyinput179);
xor g1060(G54, xenc180, keyinput180);
xor g1061(xenc181, G388, keyinput181);
xor g1062(xenc182, G1456, keyinput182);
xor g1063(xenc183, G545, keyinput183);
xnor g1064(xenc184, G893, keyinput184);
xnor g1065(xenc185, G1210, keyinput185);
xor g1066(xenc186, G1561, keyinput186);
xnor g1067(xenc187, G1921, keyinput187);
xor g1068(xenc188, G1828, keyinput188);
xnor g1069(xenc189, G65, keyinput189);
xnor g1070(xenc190, G1876, keyinput190);
xor g1071(xenc191, G1701, keyinput191);
xnor g1072(xenc192, G1393, keyinput192);
xnor g1073(xenc193, G1512, keyinput193);
xor g1074(xenc194, G572, keyinput194);
xnor g1075(xenc195, G1112, keyinput195);
xnor g1076(xenc196, G1370, keyinput196);
xor g1077(xenc197, G318, keyinput197);
xor g1078(G48, xenc198, keyinput198);
xor g1079(xenc199, G420, keyinput199);
xor g1080(xenc200, G1546, keyinput200);
xor g1081(xenc201, G1402, keyinput201);
xnor g1082(xenc202, G308, keyinput202);
xnor g1083(xenc203, G1474, keyinput203);
xnor g1084(xenc204, G37, keyinput204);
xnor g1085(xenc205, G1660, keyinput205);
xnor g1086(xenc206, G1183, keyinput206);
xor g1087(xenc207, G1165, keyinput207);
xnor g1088(xenc208, G731, keyinput208);
xnor g1089(xenc209, G1351, keyinput209);
xnor g1090(xenc210, G1424, keyinput210);
xor g1091(xenc211, G887, keyinput211);
xnor g1092(xenc212, G949, keyinput212);
xor g1093(xenc213, G360, keyinput213);
xnor g1094(xenc214, G41, keyinput214);
xnor g1095(xenc215, G1105, keyinput215);
xor g1096(xenc216, G1243, keyinput216);
xnor g1097(xenc217, G1621, keyinput217);
xnor g1098(xenc218, G366, keyinput218);
xnor g1099(xenc219, G1549, keyinput219);
xnor g1100(xenc220, G2, keyinput220);
xor g1101(G27, xenc221, keyinput221);
xnor g1102(xenc222, G268, keyinput222);
xor g1103(xenc223, G1785, keyinput223);
xor g1104(xenc224, G1466, keyinput224);
xor g1105(xenc225, G1924, keyinput225);
xor g1106(xenc226, G1216, keyinput226);
xnor g1107(xenc227, G788, keyinput227);
xnor g1108(xenc228, G1049, keyinput228);
xor g1109(xenc229, G1222, keyinput229);
xor g1110(xenc230, G1317, keyinput230);
xor g1111(xenc231, G1554, keyinput231);
xnor g1112(G21, xenc232, keyinput232);
xor g1113(xenc233, G1087, keyinput233);
xnor g1114(xenc234, G1643, keyinput234);
xor g1115(xenc235, G1533, keyinput235);
xor g1116(xenc236, G1252, keyinput236);
xnor g1117(xenc237, G1788, keyinput237);
xnor g1118(xenc238, G1437, keyinput238);
xor g1119(xenc239, G1854, keyinput239);
xnor g1120(xenc240, G58, keyinput240);
xnor g1121(xenc241, G1187, keyinput241);
xor g1122(xenc242, G984, keyinput242);
xnor g1123(xenc243, G1609, keyinput243);
xor g1124(xenc244, G198, keyinput244);
xor g1125(xenc245, G1137, keyinput245);
xor g1126(xenc246, G160, keyinput246);
xor g1127(xenc247, G1343, keyinput247);
xor g1128(xenc248, G373, keyinput248);
xor g1129(xenc249, G532, keyinput249);
xor g1130(xenc250, G1056, keyinput250);
xnor g1131(xenc251, G40, keyinput251);
xnor g1132(xenc252, G1740, keyinput252);
xor g1133(xenc253, G59, keyinput253);
xor g1134(xenc254, G943, keyinput254);
xnor g1135(xenc255, G1661, keyinput255);
endmodule
