
module c7552 ( N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, 
        N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, 
        N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, 
        N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, 
        N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, 
        N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, 
        N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, 
        N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, 
        N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, 
        N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
        N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, 
        N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, 
        N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
        N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, 
        N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, 
        N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, 
        N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, 
        N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, 
        N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, 
        N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, 
        N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, 
        N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, 
        N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, 
        N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, 
        N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, 
        N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, 
        N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, 
        N11333, N11334, N11340, N11342, N241_O, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31
 );
  input N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47,
         N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110,
         N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133,
         N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245,
         N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280,
         N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316,
         N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349,
         N352, N355, N358, N361, N364, N367, N382, N241_I, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31;
  output N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507,
         N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543,
         N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567,
         N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884,
         N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490,
         N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111,
         N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576,
         N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713,
         N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760,
         N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840,
         N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908,
         N11333, N11334, N11340, N11342, N241_O;
  wire   N1, N106, N248, N251, N254, N257, N260, N263, N267, N274, N277, N280,
         N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316,
         N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349,
         N352, N355, N358, N361, N364, N241_I, N10628, N10706, N10759, N10837,
         N10839, N582, N1113, N1112, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673;
  assign N1490 = N1;
  assign N889 = N1;
  assign N388 = N1;
  assign N387 = N1;
  assign N945 = N106;
  assign N478 = N248;
  assign N643 = N251;
  assign N482 = N254;
  assign N484 = N257;
  assign N486 = N260;
  assign N489 = N263;
  assign N492 = N267;
  assign N501 = N274;
  assign N707 = N277;
  assign N505 = N280;
  assign N507 = N283;
  assign N509 = N286;
  assign N511 = N289;
  assign N513 = N293;
  assign N515 = N296;
  assign N517 = N299;
  assign N519 = N303;
  assign N535 = N307;
  assign N537 = N310;
  assign N539 = N313;
  assign N541 = N316;
  assign N543 = N319;
  assign N545 = N322;
  assign N547 = N325;
  assign N549 = N328;
  assign N551 = N331;
  assign N553 = N334;
  assign N556 = N337;
  assign N813 = N340;
  assign N559 = N343;
  assign N561 = N346;
  assign N563 = N349;
  assign N565 = N352;
  assign N567 = N355;
  assign N569 = N358;
  assign N571 = N361;
  assign N573 = N364;
  assign N241_O = N241_I;
  assign N10102 = N10628;
  assign N10103 = N10628;
  assign N10104 = N10706;
  assign N10101 = N10759;
  assign N10838 = N10837;
  assign N10840 = N10839;
  assign N1114 = N582;
  assign N1111 = N582;
  assign N1489 = N1113;
  assign N1110 = N1112;

  OR2X1 U938 ( .IN1(N5), .IN2(N57), .Q(N881) );
  INVX0 U939 ( .INP(N15), .ZN(N582) );
  AND2X1 U940 ( .IN1(N163), .IN2(N1), .Q(N1781) );
  XOR2X1 U941 ( .IN1(n915), .IN2(n916), .Q(N11342) );
  MUX21X1 U942 ( .IN1(n917), .IN2(n918), .S(N367), .Q(n916) );
  XOR3X1 U943 ( .IN1(n919), .IN2(n920), .IN3(n921), .Q(n918) );
  XNOR2X1 U944 ( .IN1(n922), .IN2(n923), .Q(n921) );
  OA21X1 U945 ( .IN1(n924), .IN2(n925), .IN3(n926), .Q(n922) );
  MUX21X1 U946 ( .IN1(n927), .IN2(n928), .S(n929), .Q(n926) );
  NAND2X0 U947 ( .IN1(n924), .IN2(n930), .QN(n928) );
  XNOR2X1 U948 ( .IN1(n930), .IN2(n929), .Q(n925) );
  XNOR3X1 U949 ( .IN1(n931), .IN2(n932), .IN3(n933), .Q(n929) );
  XOR2X1 U950 ( .IN1(n934), .IN2(n935), .Q(n933) );
  AOI21X1 U951 ( .IN1(n924), .IN2(n936), .IN3(n937), .QN(n935) );
  NOR2X0 U952 ( .IN1(n936), .IN2(n938), .QN(n931) );
  INVX0 U953 ( .INP(n939), .ZN(n936) );
  NOR2X0 U954 ( .IN1(n940), .IN2(n941), .QN(n920) );
  XOR3X1 U955 ( .IN1(n942), .IN2(n943), .IN3(n944), .Q(n917) );
  XOR2X1 U956 ( .IN1(n938), .IN2(n945), .Q(n944) );
  NOR2X0 U957 ( .IN1(n946), .IN2(n919), .QN(n945) );
  XOR3X1 U958 ( .IN1(n947), .IN2(n930), .IN3(n948), .Q(n943) );
  XOR2X1 U959 ( .IN1(n941), .IN2(n937), .Q(n948) );
  XNOR2X1 U960 ( .IN1(n923), .IN2(n932), .Q(n942) );
  MUX21X1 U961 ( .IN1(n949), .IN2(n950), .S(n951), .Q(n915) );
  OA21X1 U962 ( .IN1(n952), .IN2(n953), .IN3(n954), .Q(n951) );
  INVX0 U963 ( .INP(n955), .ZN(n954) );
  XOR2X1 U964 ( .IN1(keyinput23), .IN2(n956), .Q(n953) );
  XOR3X1 U965 ( .IN1(n957), .IN2(n958), .IN3(n959), .Q(n950) );
  XOR2X1 U966 ( .IN1(n960), .IN2(n961), .Q(n959) );
  XOR3X1 U967 ( .IN1(n962), .IN2(n963), .IN3(n964), .Q(n958) );
  AOI21X1 U968 ( .IN1(n965), .IN2(n966), .IN3(n967), .QN(n957) );
  XOR3X1 U969 ( .IN1(n968), .IN2(n969), .IN3(n970), .Q(n949) );
  XOR2X1 U970 ( .IN1(n966), .IN2(n971), .Q(n970) );
  OA21X1 U971 ( .IN1(n972), .IN2(n964), .IN3(n973), .Q(n971) );
  XOR3X1 U972 ( .IN1(n962), .IN2(n974), .IN3(n975), .Q(n969) );
  INVX0 U973 ( .INP(n965), .ZN(n974) );
  MUX21X1 U974 ( .IN1(n961), .IN2(n972), .S(n976), .Q(n968) );
  XOR2X1 U975 ( .IN1(n977), .IN2(n978), .Q(N11340) );
  MUX21X1 U976 ( .IN1(n979), .IN2(n980), .S(n981), .Q(n978) );
  XOR2X1 U977 ( .IN1(n982), .IN2(n983), .Q(n980) );
  XOR3X1 U978 ( .IN1(n984), .IN2(n985), .IN3(n986), .Q(n983) );
  XNOR2X1 U979 ( .IN1(n987), .IN2(n988), .Q(n986) );
  NOR2X0 U980 ( .IN1(n989), .IN2(n990), .QN(n987) );
  XOR3X1 U981 ( .IN1(n991), .IN2(n992), .IN3(n993), .Q(n982) );
  XNOR2X1 U982 ( .IN1(n994), .IN2(n995), .Q(n993) );
  AOI21X1 U983 ( .IN1(n988), .IN2(n996), .IN3(n997), .QN(n994) );
  NOR2X0 U984 ( .IN1(n996), .IN2(n998), .QN(n992) );
  INVX0 U985 ( .INP(n999), .ZN(n996) );
  XOR2X1 U986 ( .IN1(n1000), .IN2(n1001), .Q(n979) );
  XNOR3X1 U987 ( .IN1(n988), .IN2(n1002), .IN3(n997), .Q(n1001) );
  AO21X1 U988 ( .IN1(n988), .IN2(n998), .IN3(n1003), .Q(n997) );
  XOR2X1 U989 ( .IN1(n984), .IN2(n985), .Q(n1002) );
  XOR2X1 U990 ( .IN1(n1004), .IN2(n1005), .Q(n985) );
  XOR3X1 U991 ( .IN1(n1006), .IN2(n990), .IN3(n1007), .Q(n1000) );
  XOR2X1 U992 ( .IN1(n998), .IN2(n991), .Q(n1007) );
  MUX21X1 U993 ( .IN1(n1008), .IN2(n1009), .S(n1010), .Q(n977) );
  NOR2X0 U994 ( .IN1(n1011), .IN2(n1012), .QN(n1010) );
  AND3X1 U995 ( .IN1(n1013), .IN2(n981), .IN3(n988), .Q(n1011) );
  XOR3X1 U996 ( .IN1(n1014), .IN2(n1015), .IN3(n1016), .Q(n1009) );
  XOR3X1 U997 ( .IN1(n1017), .IN2(n1018), .IN3(n1019), .Q(n1016) );
  XOR3X1 U998 ( .IN1(n1020), .IN2(n1014), .IN3(n1021), .Q(n1008) );
  XNOR3X1 U999 ( .IN1(keyinput28), .IN2(n1015), .IN3(n1022), .Q(n1021) );
  AO21X1 U1000 ( .IN1(n1023), .IN2(n1024), .IN3(n1025), .Q(n1015) );
  XOR2X1 U1001 ( .IN1(n1026), .IN2(n1027), .Q(n1014) );
  MUX21X1 U1002 ( .IN1(n1028), .IN2(n1029), .S(n1030), .Q(n1020) );
  XOR2X1 U1003 ( .IN1(n1031), .IN2(n1032), .Q(N11334) );
  MUX21X1 U1004 ( .IN1(n1033), .IN2(n1034), .S(n1035), .Q(n1032) );
  XOR2X1 U1005 ( .IN1(n1036), .IN2(n1037), .Q(n1034) );
  XNOR3X1 U1006 ( .IN1(n1038), .IN2(n1039), .IN3(n1040), .Q(n1037) );
  NOR2X0 U1007 ( .IN1(n1041), .IN2(n1042), .QN(n1038) );
  XOR3X1 U1008 ( .IN1(n1043), .IN2(n1044), .IN3(n1045), .Q(n1036) );
  XOR2X1 U1009 ( .IN1(n1046), .IN2(n1047), .Q(n1045) );
  NOR2X0 U1010 ( .IN1(n1048), .IN2(n1049), .QN(n1047) );
  NAND3X0 U1011 ( .IN1(n1050), .IN2(n1051), .IN3(n1052), .QN(n1046) );
  NAND2X0 U1012 ( .IN1(n1053), .IN2(n1054), .QN(n1051) );
  XNOR2X1 U1013 ( .IN1(keyinput13), .IN2(n1055), .Q(n1050) );
  NAND2X0 U1014 ( .IN1(n1056), .IN2(n1057), .QN(n1043) );
  XOR2X1 U1015 ( .IN1(n1058), .IN2(n1059), .Q(n1033) );
  XOR3X1 U1016 ( .IN1(n1039), .IN2(n1040), .IN3(n1060), .Q(n1059) );
  XOR2X1 U1017 ( .IN1(n1061), .IN2(n1062), .Q(n1060) );
  NAND2X0 U1018 ( .IN1(keyinput29), .IN2(n1042), .QN(n1062) );
  XOR2X1 U1019 ( .IN1(n1063), .IN2(n1064), .Q(n1040) );
  XOR3X1 U1020 ( .IN1(n1065), .IN2(n1066), .IN3(n1067), .Q(n1058) );
  XOR2X1 U1021 ( .IN1(n1068), .IN2(n1054), .Q(n1066) );
  MUX21X1 U1022 ( .IN1(n1069), .IN2(n1070), .S(n1071), .Q(n1031) );
  XOR2X1 U1023 ( .IN1(n1072), .IN2(n1073), .Q(n1070) );
  XOR2X1 U1024 ( .IN1(n1072), .IN2(n1074), .Q(n1069) );
  XNOR2X1 U1025 ( .IN1(n1075), .IN2(n1076), .Q(n1072) );
  XOR2X1 U1026 ( .IN1(n1077), .IN2(n1078), .Q(N11333) );
  MUX21X1 U1027 ( .IN1(n1079), .IN2(n1080), .S(n1081), .Q(n1078) );
  XOR3X1 U1028 ( .IN1(n1082), .IN2(n1083), .IN3(n1084), .Q(n1080) );
  XOR3X1 U1029 ( .IN1(n1085), .IN2(n1086), .IN3(n1087), .Q(n1084) );
  XNOR3X1 U1030 ( .IN1(n1088), .IN2(n1089), .IN3(n1090), .Q(n1087) );
  NOR2X0 U1031 ( .IN1(n1091), .IN2(n1092), .QN(n1089) );
  XOR3X1 U1032 ( .IN1(n1093), .IN2(n1094), .IN3(n1095), .Q(n1085) );
  AOI21X1 U1033 ( .IN1(n1082), .IN2(n1091), .IN3(n1096), .QN(n1095) );
  AOI21X1 U1034 ( .IN1(n1097), .IN2(n1091), .IN3(n1098), .QN(n1083) );
  XOR3X1 U1035 ( .IN1(n1099), .IN2(n1100), .IN3(n1101), .Q(n1079) );
  XNOR3X1 U1036 ( .IN1(n1098), .IN2(n1092), .IN3(n1102), .Q(n1101) );
  XNOR2X1 U1037 ( .IN1(n1090), .IN2(n1103), .Q(n1102) );
  NOR2X0 U1038 ( .IN1(n1104), .IN2(n1093), .QN(n1103) );
  XOR2X1 U1039 ( .IN1(n1096), .IN2(n1105), .Q(n1100) );
  XOR2X1 U1040 ( .IN1(n1082), .IN2(n1094), .Q(n1099) );
  OA21X1 U1041 ( .IN1(n1106), .IN2(n1107), .IN3(n1108), .Q(n1077) );
  MUX21X1 U1042 ( .IN1(n1109), .IN2(n1110), .S(n1111), .Q(n1108) );
  NAND2X0 U1043 ( .IN1(n1112), .IN2(n1113), .QN(n1110) );
  XOR2X1 U1044 ( .IN1(keyinput19), .IN2(n1114), .Q(n1113) );
  NAND2X0 U1045 ( .IN1(n1115), .IN2(n1107), .QN(n1109) );
  MUX21X1 U1046 ( .IN1(n1115), .IN2(n1112), .S(n1111), .Q(n1106) );
  XOR3X1 U1047 ( .IN1(n1116), .IN2(n1117), .IN3(n1118), .Q(n1112) );
  XOR3X1 U1048 ( .IN1(keyinput31), .IN2(n1119), .IN3(n1120), .Q(n1117) );
  OA21X1 U1049 ( .IN1(n1121), .IN2(n1122), .IN3(n1123), .Q(n1120) );
  XOR2X1 U1050 ( .IN1(n1124), .IN2(keyinput22), .Q(n1123) );
  NAND2X0 U1051 ( .IN1(n1122), .IN2(n1121), .QN(n1124) );
  XOR2X1 U1052 ( .IN1(n1125), .IN2(n1126), .Q(n1115) );
  XOR3X1 U1053 ( .IN1(n1119), .IN2(n1127), .IN3(n1128), .Q(n1126) );
  XOR2X1 U1054 ( .IN1(n1129), .IN2(n1130), .Q(n1125) );
  NAND3X0 U1055 ( .IN1(N133), .IN2(n1131), .IN3(N134), .QN(N1113) );
  NAND2X0 U1056 ( .IN1(N242), .IN2(n1131), .QN(N1112) );
  INVX0 U1057 ( .INP(N5), .ZN(n1131) );
  XNOR2X1 U1058 ( .IN1(n1024), .IN2(n1132), .Q(N10908) );
  XOR2X1 U1059 ( .IN1(n1023), .IN2(n1133), .Q(N10907) );
  AOI21X1 U1060 ( .IN1(n1030), .IN2(n1132), .IN3(n1017), .QN(n1133) );
  MUX21X1 U1061 ( .IN1(n1134), .IN2(n1135), .S(n1132), .Q(N10906) );
  AO21X1 U1062 ( .IN1(n1136), .IN2(n1137), .IN3(n1138), .Q(n1135) );
  XOR2X1 U1063 ( .IN1(n1139), .IN2(keyinput24), .Q(n1138) );
  NAND2X0 U1064 ( .IN1(n1029), .IN2(n1027), .QN(n1139) );
  INVX0 U1065 ( .INP(n1029), .ZN(n1136) );
  NOR2X0 U1066 ( .IN1(n1028), .IN2(n1025), .QN(n1029) );
  XOR2X1 U1067 ( .IN1(n1137), .IN2(n1018), .Q(n1134) );
  INVX0 U1068 ( .INP(n1028), .ZN(n1018) );
  XOR2X1 U1069 ( .IN1(n1140), .IN2(n1141), .Q(N10905) );
  OA21X1 U1070 ( .IN1(n1019), .IN2(n1132), .IN3(n1022), .Q(n1141) );
  NAND2X0 U1071 ( .IN1(n1142), .IN2(n1143), .QN(n1022) );
  INVX0 U1072 ( .INP(n1019), .ZN(n1142) );
  NAND2X0 U1073 ( .IN1(n1144), .IN2(n1145), .QN(n1132) );
  NAND3X0 U1074 ( .IN1(n984), .IN2(n1146), .IN3(n1147), .QN(n1145) );
  XOR2X1 U1075 ( .IN1(n1148), .IN2(n1004), .Q(N10871) );
  NAND2X0 U1076 ( .IN1(n1006), .IN2(n1149), .QN(n1148) );
  MUX21X1 U1077 ( .IN1(n1150), .IN2(n1151), .S(keyinput30), .Q(N10870) );
  XOR2X1 U1078 ( .IN1(n1152), .IN2(n1153), .Q(n1151) );
  AO21X1 U1079 ( .IN1(n1153), .IN2(n1152), .IN3(n1154), .Q(n1150) );
  XOR2X1 U1080 ( .IN1(n1146), .IN2(n1155), .Q(N10869) );
  OR2X1 U1081 ( .IN1(n998), .IN2(n1147), .Q(n1155) );
  AND2X1 U1082 ( .IN1(n1156), .IN2(n1005), .Q(n1147) );
  XOR2X1 U1083 ( .IN1(n1157), .IN2(n1158), .Q(N10868) );
  NOR2X0 U1084 ( .IN1(n1003), .IN2(n1159), .QN(n1158) );
  OA21X1 U1085 ( .IN1(n1160), .IN2(n1154), .IN3(n1146), .Q(n1159) );
  NOR2X0 U1086 ( .IN1(n1152), .IN2(n1153), .QN(n1154) );
  NOR2X0 U1087 ( .IN1(n990), .IN2(n1156), .QN(n1153) );
  NOR2X0 U1088 ( .IN1(n1149), .IN2(n1161), .QN(n1156) );
  NAND2X0 U1089 ( .IN1(n991), .IN2(n1162), .QN(n1149) );
  XOR2X1 U1090 ( .IN1(n1162), .IN2(n991), .Q(N10827) );
  XOR2X1 U1091 ( .IN1(n1163), .IN2(n1076), .Q(N10839) );
  XNOR2X1 U1092 ( .IN1(n1164), .IN2(n1165), .Q(N10837) );
  OA21X1 U1093 ( .IN1(n1074), .IN2(n1163), .IN3(n1166), .Q(n1165) );
  INVX0 U1094 ( .INP(n1073), .ZN(n1166) );
  XOR2X1 U1095 ( .IN1(n1167), .IN2(n1119), .Q(N10763) );
  MUX21X1 U1096 ( .IN1(n1130), .IN2(n1168), .S(n1167), .Q(N10762) );
  XOR2X1 U1097 ( .IN1(n1122), .IN2(n1116), .Q(n1168) );
  XOR2X1 U1098 ( .IN1(n1116), .IN2(n1169), .Q(n1130) );
  XOR2X1 U1099 ( .IN1(n1114), .IN2(n1170), .Q(N10761) );
  OA21X1 U1100 ( .IN1(n1128), .IN2(n1167), .IN3(n1121), .Q(n1170) );
  AO21X1 U1101 ( .IN1(n1119), .IN2(n1116), .IN3(n1128), .Q(n1121) );
  MUX21X1 U1102 ( .IN1(n1171), .IN2(n1118), .S(n1167), .Q(N10760) );
  XOR2X1 U1103 ( .IN1(n1127), .IN2(n1172), .Q(n1118) );
  NOR2X0 U1104 ( .IN1(n1173), .IN2(n1174), .QN(n1172) );
  XOR2X1 U1105 ( .IN1(n1174), .IN2(n1175), .Q(n1171) );
  AO221X1 U1106 ( .IN1(n1176), .IN2(n1076), .IN3(N38), .IN4(n1177), .IN5(n1074), .Q(N10759) );
  NOR2X0 U1107 ( .IN1(n1178), .IN2(n1164), .QN(n1176) );
  INVX0 U1108 ( .INP(n1163), .ZN(n1178) );
  AO21X1 U1109 ( .IN1(n1179), .IN2(n1039), .IN3(n1180), .Q(n1163) );
  OR4X1 U1110 ( .IN1(N10575), .IN2(N10576), .IN3(N10574), .IN4(n1181), .Q(
        N10729) );
  OR4X1 U1111 ( .IN1(N885), .IN2(N884), .IN3(N883), .IN4(N882), .Q(n1181) );
  NAND4X0 U1112 ( .IN1(N240), .IN2(N228), .IN3(N184), .IN4(N150), .QN(N882) );
  NAND4X0 U1113 ( .IN1(N230), .IN2(N218), .IN3(N210), .IN4(N152), .QN(N883) );
  NAND4X0 U1114 ( .IN1(N186), .IN2(N185), .IN3(N183), .IN4(N182), .QN(N884) );
  NAND4X0 U1115 ( .IN1(N199), .IN2(N188), .IN3(N172), .IN4(N162), .QN(N885) );
  XOR2X1 U1116 ( .IN1(n1182), .IN2(n1183), .Q(N10718) );
  NAND2X0 U1117 ( .IN1(n1184), .IN2(n1185), .QN(n1182) );
  MUX21X1 U1118 ( .IN1(n1186), .IN2(n1187), .S(n1188), .Q(N10717) );
  OA21X1 U1119 ( .IN1(n1064), .IN2(n1185), .IN3(n1065), .Q(n1187) );
  INVX0 U1120 ( .INP(n1049), .ZN(n1065) );
  NAND2X0 U1121 ( .IN1(n1042), .IN2(n1189), .QN(n1185) );
  AO21X1 U1122 ( .IN1(n1048), .IN2(n1189), .IN3(n1049), .Q(n1186) );
  XOR2X1 U1123 ( .IN1(n1190), .IN2(n1054), .Q(N10716) );
  NAND2X0 U1124 ( .IN1(n1056), .IN2(n1191), .QN(n1190) );
  INVX0 U1125 ( .INP(n1067), .ZN(n1056) );
  XNOR2X1 U1126 ( .IN1(n1039), .IN2(n1192), .Q(N10715) );
  NOR2X0 U1127 ( .IN1(n1179), .IN2(n1061), .QN(n1192) );
  NAND2X0 U1128 ( .IN1(n1052), .IN2(n1055), .QN(n1061) );
  NAND4X0 U1129 ( .IN1(n1054), .IN2(n1188), .IN3(n1068), .IN4(n1183), .QN(
        n1055) );
  AOI21X1 U1130 ( .IN1(n1054), .IN2(n1193), .IN3(n1194), .QN(n1052) );
  AO21X1 U1131 ( .IN1(n1195), .IN2(n1188), .IN3(n1196), .Q(n1193) );
  NOR2X0 U1132 ( .IN1(n1191), .IN2(n1044), .QN(n1179) );
  NAND2X0 U1133 ( .IN1(n1053), .IN2(n1189), .QN(n1191) );
  XOR2X1 U1134 ( .IN1(n1086), .IN2(n1197), .Q(N10714) );
  NOR2X0 U1135 ( .IN1(n1198), .IN2(keyinput17), .QN(n1197) );
  AOI21X1 U1136 ( .IN1(n1199), .IN2(n1093), .IN3(n1104), .QN(n1198) );
  XOR2X1 U1137 ( .IN1(n1200), .IN2(n1082), .Q(N10713) );
  OR2X1 U1138 ( .IN1(n1092), .IN2(n1201), .Q(n1200) );
  XOR2X1 U1139 ( .IN1(n1202), .IN2(n1203), .Q(N10712) );
  AOI21X1 U1140 ( .IN1(n1082), .IN2(n1201), .IN3(n1096), .QN(n1203) );
  NAND3X0 U1141 ( .IN1(n1204), .IN2(n1205), .IN3(n1206), .QN(n1096) );
  NAND2X0 U1142 ( .IN1(n1207), .IN2(n1082), .QN(n1206) );
  INVX0 U1143 ( .INP(n1208), .ZN(n1201) );
  XNOR2X1 U1144 ( .IN1(n1090), .IN2(n1209), .Q(N10711) );
  NOR2X0 U1145 ( .IN1(n1210), .IN2(n1098), .QN(n1209) );
  AO221X1 U1146 ( .IN1(n1207), .IN2(n1097), .IN3(n1211), .IN4(n1094), .IN5(
        n1212), .Q(n1098) );
  INVX0 U1147 ( .INP(n1204), .ZN(n1211) );
  NAND3X0 U1148 ( .IN1(n1086), .IN2(n1082), .IN3(n1104), .QN(n1204) );
  AO22X1 U1149 ( .IN1(N38), .IN2(n1177), .IN3(n1075), .IN4(n1213), .Q(N10706)
         );
  AO21X1 U1150 ( .IN1(n1076), .IN2(n1071), .IN3(n1074), .Q(n1213) );
  OR2X1 U1151 ( .IN1(n1180), .IN2(n1214), .Q(n1071) );
  AND4X1 U1152 ( .IN1(n1053), .IN2(n1054), .IN3(n1039), .IN4(n1035), .Q(n1214)
         );
  NAND2X0 U1153 ( .IN1(n1215), .IN2(n1216), .QN(n1035) );
  NAND3X0 U1154 ( .IN1(n1175), .IN2(n1111), .IN3(n1173), .QN(n1216) );
  OR2X1 U1155 ( .IN1(n1217), .IN2(n1218), .Q(n1111) );
  AND4X1 U1156 ( .IN1(n1091), .IN2(n1097), .IN3(n1090), .IN4(n1081), .Q(n1218)
         );
  AO21X1 U1157 ( .IN1(n1219), .IN2(n1220), .IN3(n1221), .Q(n1081) );
  NAND2X0 U1158 ( .IN1(n1222), .IN2(n1223), .QN(n1220) );
  NAND3X0 U1159 ( .IN1(n988), .IN2(n981), .IN3(n1013), .QN(n1223) );
  AO21X1 U1160 ( .IN1(n962), .IN2(n1224), .IN3(n1225), .Q(n981) );
  INVX0 U1161 ( .INP(n1226), .ZN(n1225) );
  NAND2X0 U1162 ( .IN1(n960), .IN2(n1227), .QN(n1224) );
  NAND3X0 U1163 ( .IN1(n975), .IN2(n1228), .IN3(n967), .QN(n1227) );
  OA21X1 U1164 ( .IN1(n964), .IN2(n1229), .IN3(n973), .Q(n960) );
  INVX0 U1165 ( .INP(n975), .ZN(n964) );
  OA21X1 U1166 ( .IN1(n1230), .IN2(n1231), .IN3(n973), .Q(n975) );
  INVX0 U1167 ( .INP(n1012), .ZN(n1222) );
  NAND2X0 U1168 ( .IN1(n1232), .IN2(n1233), .QN(n1012) );
  NAND3X0 U1169 ( .IN1(n984), .IN2(n998), .IN3(n988), .QN(n1233) );
  XOR2X1 U1170 ( .IN1(N349), .IN2(n1234), .Q(n988) );
  INVX0 U1171 ( .INP(n1057), .ZN(n1053) );
  NAND2X0 U1172 ( .IN1(n1048), .IN2(n1188), .QN(n1057) );
  AND2X1 U1173 ( .IN1(n1042), .IN2(n1183), .Q(n1048) );
  AO22X1 U1174 ( .IN1(n1235), .IN2(n1236), .IN3(n1039), .IN4(n1237), .Q(n1180)
         );
  AO21X1 U1175 ( .IN1(n1054), .IN2(n1067), .IN3(n1194), .Q(n1237) );
  AO21X1 U1176 ( .IN1(n1188), .IN2(n1049), .IN3(n1196), .Q(n1067) );
  AO21X1 U1177 ( .IN1(n1068), .IN2(n1183), .IN3(n1195), .Q(n1049) );
  INVX0 U1178 ( .INP(n1064), .ZN(n1183) );
  AO21X1 U1179 ( .IN1(N254), .IN2(n1238), .IN3(n1195), .Q(n1064) );
  NOR2X0 U1180 ( .IN1(n1238), .IN2(N254), .QN(n1195) );
  INVX0 U1181 ( .INP(n1063), .ZN(n1188) );
  AO21X1 U1182 ( .IN1(N106), .IN2(n1239), .IN3(n1196), .Q(n1063) );
  NOR2X0 U1183 ( .IN1(N106), .IN2(n1239), .QN(n1196) );
  INVX0 U1184 ( .INP(n1044), .ZN(n1054) );
  AO21X1 U1185 ( .IN1(N257), .IN2(n1240), .IN3(n1194), .Q(n1044) );
  NOR2X0 U1186 ( .IN1(n1240), .IN2(N257), .QN(n1194) );
  XOR2X1 U1187 ( .IN1(n1236), .IN2(n1235), .Q(n1039) );
  NOR2X0 U1188 ( .IN1(n1074), .IN2(n1073), .QN(n1076) );
  NOR3X0 U1189 ( .IN1(n1241), .IN2(N38), .IN3(n1242), .QN(n1073) );
  OA21X1 U1190 ( .IN1(n1242), .IN2(n1241), .IN3(N38), .Q(n1074) );
  XOR2X1 U1191 ( .IN1(n1164), .IN2(keyinput3), .Q(n1075) );
  XNOR2X1 U1192 ( .IN1(n1177), .IN2(N38), .Q(n1164) );
  NAND2X0 U1193 ( .IN1(N267), .IN2(N382), .QN(n1177) );
  AO21X1 U1194 ( .IN1(n1243), .IN2(n1244), .IN3(n1245), .Q(N10704) );
  INVX0 U1195 ( .INP(n1246), .ZN(n1244) );
  MUX21X1 U1196 ( .IN1(n1247), .IN2(n1248), .S(keyinput27), .Q(n1243) );
  NAND2X0 U1197 ( .IN1(n1249), .IN2(n1250), .QN(n1248) );
  INVX0 U1198 ( .INP(n1251), .ZN(n1249) );
  INVX0 U1199 ( .INP(n1252), .ZN(n1247) );
  XOR2X1 U1200 ( .IN1(n1189), .IN2(n1042), .Q(N10641) );
  NOR2X0 U1201 ( .IN1(n1068), .IN2(n1041), .QN(n1042) );
  NOR2X0 U1202 ( .IN1(n1253), .IN2(n1254), .QN(n1041) );
  INVX0 U1203 ( .INP(n1184), .ZN(n1068) );
  NAND2X0 U1204 ( .IN1(n1254), .IN2(n1253), .QN(n1184) );
  NAND2X0 U1205 ( .IN1(n1215), .IN2(n1255), .QN(n1189) );
  NAND3X0 U1206 ( .IN1(n1175), .IN2(n1167), .IN3(n1173), .QN(n1255) );
  AND3X1 U1207 ( .IN1(n1116), .IN2(n1114), .IN3(n1119), .Q(n1173) );
  NOR2X0 U1208 ( .IN1(n1169), .IN2(n1256), .QN(n1119) );
  INVX0 U1209 ( .INP(n1122), .ZN(n1256) );
  NAND2X0 U1210 ( .IN1(N293), .IN2(n1257), .QN(n1122) );
  AO21X1 U1211 ( .IN1(n1210), .IN2(n1090), .IN3(n1217), .Q(n1167) );
  AO22X1 U1212 ( .IN1(n1258), .IN2(n1259), .IN3(n1090), .IN4(n1260), .Q(n1217)
         );
  AO21X1 U1213 ( .IN1(n1097), .IN2(n1092), .IN3(n1212), .Q(n1260) );
  AO21X1 U1214 ( .IN1(n1094), .IN2(n1261), .IN3(n1262), .Q(n1212) );
  INVX0 U1215 ( .INP(n1205), .ZN(n1261) );
  AO21X1 U1216 ( .IN1(n1104), .IN2(n1086), .IN3(n1207), .Q(n1092) );
  INVX0 U1217 ( .INP(n1263), .ZN(n1097) );
  XOR2X1 U1218 ( .IN1(n1259), .IN2(n1258), .Q(n1090) );
  NOR2X0 U1219 ( .IN1(n1208), .IN2(n1263), .QN(n1210) );
  NAND2X0 U1220 ( .IN1(n1082), .IN2(n1094), .QN(n1263) );
  INVX0 U1221 ( .INP(n1202), .ZN(n1094) );
  AO21X1 U1222 ( .IN1(N286), .IN2(n1264), .IN3(n1262), .Q(n1202) );
  NOR2X0 U1223 ( .IN1(n1264), .IN2(N286), .QN(n1262) );
  INVX0 U1224 ( .INP(n1265), .ZN(n1264) );
  OA21X1 U1225 ( .IN1(n1266), .IN2(n1267), .IN3(n1205), .Q(n1082) );
  NAND2X0 U1226 ( .IN1(n1267), .IN2(n1266), .QN(n1205) );
  NAND2X0 U1227 ( .IN1(n1091), .IN2(n1199), .QN(n1208) );
  AND2X1 U1228 ( .IN1(n1093), .IN2(n1086), .Q(n1091) );
  INVX0 U1229 ( .INP(n1105), .ZN(n1086) );
  AO21X1 U1230 ( .IN1(N280), .IN2(n1268), .IN3(n1207), .Q(n1105) );
  NOR2X0 U1231 ( .IN1(n1268), .IN2(N280), .QN(n1207) );
  INVX0 U1232 ( .INP(n1269), .ZN(n1268) );
  OA22X1 U1233 ( .IN1(n1270), .IN2(N303), .IN3(n1127), .IN4(n1129), .Q(n1215)
         );
  INVX0 U1234 ( .INP(n1174), .ZN(n1129) );
  AO21X1 U1235 ( .IN1(n1114), .IN2(n1128), .IN3(n1271), .Q(n1174) );
  AO22X1 U1236 ( .IN1(n1272), .IN2(n1273), .IN3(n1169), .IN4(n1116), .Q(n1128)
         );
  XOR2X1 U1237 ( .IN1(n1273), .IN2(n1272), .Q(n1116) );
  NOR2X0 U1238 ( .IN1(n1257), .IN2(N293), .QN(n1169) );
  INVX0 U1239 ( .INP(n1274), .ZN(n1257) );
  INVX0 U1240 ( .INP(n1107), .ZN(n1114) );
  AO21X1 U1241 ( .IN1(N299), .IN2(n1275), .IN3(n1271), .Q(n1107) );
  NOR2X0 U1242 ( .IN1(N299), .IN2(n1275), .QN(n1271) );
  INVX0 U1243 ( .INP(n1175), .ZN(n1127) );
  XOR2X1 U1244 ( .IN1(N303), .IN2(n1270), .Q(n1175) );
  XOR2X1 U1245 ( .IN1(n1199), .IN2(n1093), .Q(N10632) );
  NOR2X0 U1246 ( .IN1(n1088), .IN2(n1104), .QN(n1093) );
  AND2X1 U1247 ( .IN1(n1276), .IN2(n1277), .Q(n1104) );
  NOR2X0 U1248 ( .IN1(n1277), .IN2(n1276), .QN(n1088) );
  AO21X1 U1249 ( .IN1(n1219), .IN2(n1278), .IN3(n1221), .Q(n1199) );
  AO21X1 U1250 ( .IN1(n1140), .IN2(n1019), .IN3(n1279), .Q(n1221) );
  AO21X1 U1251 ( .IN1(n1027), .IN2(n1028), .IN3(n1280), .Q(n1019) );
  AO22X1 U1252 ( .IN1(n1281), .IN2(n1282), .IN3(n1017), .IN4(n1283), .Q(n1028)
         );
  INVX0 U1253 ( .INP(n1023), .ZN(n1283) );
  INVX0 U1254 ( .INP(n1026), .ZN(n1140) );
  NAND2X0 U1255 ( .IN1(n1144), .IN2(n1284), .QN(n1278) );
  NAND3X0 U1256 ( .IN1(n1162), .IN2(n1146), .IN3(n1013), .QN(n1284) );
  NOR2X0 U1257 ( .IN1(n999), .IN2(n1157), .QN(n1013) );
  NAND2X0 U1258 ( .IN1(n989), .IN2(n1005), .QN(n999) );
  AND2X1 U1259 ( .IN1(n991), .IN2(n1004), .Q(n989) );
  AND2X1 U1260 ( .IN1(n1006), .IN2(n995), .Q(n991) );
  NAND2X0 U1261 ( .IN1(N340), .IN2(n1285), .QN(n995) );
  INVX0 U1262 ( .INP(n1286), .ZN(n1006) );
  NAND3X0 U1263 ( .IN1(n1287), .IN2(n1226), .IN3(n1288), .QN(n1162) );
  NAND4X0 U1264 ( .IN1(n1289), .IN2(n967), .IN3(n962), .IN4(n1228), .QN(n1288)
         );
  INVX0 U1265 ( .INP(n1290), .ZN(n1289) );
  INVX0 U1266 ( .INP(n1291), .ZN(n1287) );
  AND2X1 U1267 ( .IN1(n1232), .IN2(n1292), .Q(n1144) );
  NAND3X0 U1268 ( .IN1(n998), .IN2(n1146), .IN3(n984), .QN(n1292) );
  AO21X1 U1269 ( .IN1(N349), .IN2(n1293), .IN3(n1294), .Q(n1146) );
  XOR2X1 U1270 ( .IN1(keyinput12), .IN2(n1295), .Q(n1294) );
  NOR2X0 U1271 ( .IN1(N349), .IN2(n1293), .QN(n1295) );
  AO21X1 U1272 ( .IN1(n1005), .IN2(n990), .IN3(n1160), .Q(n998) );
  AO21X1 U1273 ( .IN1(n1286), .IN2(n1004), .IN3(n1296), .Q(n990) );
  INVX0 U1274 ( .INP(n1161), .ZN(n1004) );
  AO21X1 U1275 ( .IN1(N343), .IN2(n1297), .IN3(n1296), .Q(n1161) );
  NOR2X0 U1276 ( .IN1(n1297), .IN2(N343), .QN(n1296) );
  INVX0 U1277 ( .INP(n1298), .ZN(n1297) );
  NOR2X0 U1278 ( .IN1(n1285), .IN2(N340), .QN(n1286) );
  INVX0 U1279 ( .INP(n1299), .ZN(n1285) );
  INVX0 U1280 ( .INP(n1152), .ZN(n1005) );
  AO21X1 U1281 ( .IN1(N346), .IN2(n1300), .IN3(n1160), .Q(n1152) );
  NOR2X0 U1282 ( .IN1(n1300), .IN2(N346), .QN(n1160) );
  AOI22X1 U1283 ( .IN1(n1301), .IN2(n1302), .IN3(n1003), .IN4(n984), .QN(n1232) );
  INVX0 U1284 ( .INP(n1157), .ZN(n984) );
  XOR2X1 U1285 ( .IN1(n1301), .IN2(N352), .Q(n1157) );
  NOR2X0 U1286 ( .IN1(n1234), .IN2(N349), .QN(n1003) );
  NOR2X0 U1287 ( .IN1(n1143), .IN2(n1026), .QN(n1219) );
  AO21X1 U1288 ( .IN1(N364), .IN2(n1303), .IN3(n1279), .Q(n1026) );
  NOR2X0 U1289 ( .IN1(n1303), .IN2(N364), .QN(n1279) );
  INVX0 U1290 ( .INP(n1304), .ZN(n1303) );
  NAND2X0 U1291 ( .IN1(n1025), .IN2(n1027), .QN(n1143) );
  INVX0 U1292 ( .INP(n1137), .ZN(n1027) );
  AO21X1 U1293 ( .IN1(N361), .IN2(n1305), .IN3(n1280), .Q(n1137) );
  NOR2X0 U1294 ( .IN1(n1305), .IN2(N361), .QN(n1280) );
  INVX0 U1295 ( .INP(n1306), .ZN(n1305) );
  NOR2X0 U1296 ( .IN1(n1024), .IN2(n1023), .QN(n1025) );
  XOR2X1 U1297 ( .IN1(n1281), .IN2(N358), .Q(n1023) );
  NAND2X0 U1298 ( .IN1(n1030), .IN2(n1307), .QN(n1024) );
  INVX0 U1299 ( .INP(n1017), .ZN(n1307) );
  NOR2X0 U1300 ( .IN1(n1308), .IN2(N355), .QN(n1017) );
  NAND2X0 U1301 ( .IN1(N355), .IN2(n1308), .QN(n1030) );
  INVX0 U1302 ( .INP(n1309), .ZN(n1308) );
  AO22X1 U1303 ( .IN1(N38), .IN2(n1310), .IN3(n1311), .IN4(n1312), .Q(N10628)
         );
  AO21X1 U1304 ( .IN1(N271), .IN2(N245), .IN3(n1242), .Q(n1311) );
  OR4X1 U1305 ( .IN1(n1312), .IN2(n1242), .IN3(N245), .IN4(N271), .Q(n1310) );
  INVX0 U1306 ( .INP(N382), .ZN(n1242) );
  AO221X1 U1307 ( .IN1(n1313), .IN2(n1314), .IN3(n1315), .IN4(n1316), .IN5(
        n1317), .Q(n1312) );
  OA221X1 U1308 ( .IN1(n1318), .IN2(n1319), .IN3(n1320), .IN4(n1321), .IN5(
        n1322), .Q(n1317) );
  INVX0 U1309 ( .INP(n1323), .ZN(n1322) );
  AND2X1 U1310 ( .IN1(n1318), .IN2(n1319), .Q(n1320) );
  AOI22X1 U1311 ( .IN1(n1324), .IN2(n1325), .IN3(n1326), .IN4(n1327), .QN(
        n1319) );
  OR2X1 U1312 ( .IN1(n1324), .IN2(n1325), .Q(n1327) );
  INVX0 U1313 ( .INP(n1328), .ZN(n1325) );
  AO22X1 U1314 ( .IN1(n1329), .IN2(n1330), .IN3(n1331), .IN4(n1332), .Q(n1324)
         );
  OR2X1 U1315 ( .IN1(n1329), .IN2(n1330), .Q(n1332) );
  INVX0 U1316 ( .INP(n1333), .ZN(n1330) );
  NAND2X0 U1317 ( .IN1(n1334), .IN2(n1335), .QN(n1329) );
  OA221X1 U1318 ( .IN1(n1318), .IN2(n1321), .IN3(n1336), .IN4(n1337), .IN5(
        n1338), .Q(n1314) );
  NOR2X0 U1319 ( .IN1(n1323), .IN2(n1339), .QN(n1338) );
  OA21X1 U1320 ( .IN1(n1340), .IN2(n1341), .IN3(n1342), .Q(n1339) );
  NOR2X0 U1321 ( .IN1(n1343), .IN2(n1315), .QN(n1323) );
  XOR2X1 U1322 ( .IN1(n1316), .IN2(keyinput8), .Q(n1343) );
  INVX0 U1323 ( .INP(n1341), .ZN(n1336) );
  AO22X1 U1324 ( .IN1(n1344), .IN2(n1345), .IN3(n1346), .IN4(n1347), .Q(n1341)
         );
  NAND2X0 U1325 ( .IN1(n1348), .IN2(n1349), .QN(n1347) );
  INVX0 U1326 ( .INP(n1349), .ZN(n1344) );
  AO221X1 U1327 ( .IN1(n1350), .IN2(n1351), .IN3(n1352), .IN4(n1353), .IN5(
        n1354), .Q(n1349) );
  OA221X1 U1328 ( .IN1(n1355), .IN2(n1356), .IN3(n1357), .IN4(n1358), .IN5(
        n1359), .Q(n1354) );
  AND2X1 U1329 ( .IN1(n1355), .IN2(n1356), .Q(n1357) );
  OA22X1 U1330 ( .IN1(n1360), .IN2(n1361), .IN3(n1362), .IN4(n1363), .Q(n1356)
         );
  AND2X1 U1331 ( .IN1(n1360), .IN2(n1361), .Q(n1363) );
  OA22X1 U1332 ( .IN1(n1364), .IN2(n1365), .IN3(n1366), .IN4(n1367), .Q(n1360)
         );
  AND2X1 U1333 ( .IN1(n1365), .IN2(n1364), .Q(n1367) );
  OA22X1 U1334 ( .IN1(n1368), .IN2(n1369), .IN3(n1370), .IN4(n1371), .Q(n1365)
         );
  AND2X1 U1335 ( .IN1(n1369), .IN2(n1368), .Q(n1371) );
  OA21X1 U1336 ( .IN1(n1372), .IN2(n1373), .IN3(n1374), .Q(n1369) );
  AO22X1 U1337 ( .IN1(n1372), .IN2(n1373), .IN3(n1375), .IN4(n1376), .Q(n1374)
         );
  OA221X1 U1338 ( .IN1(n1364), .IN2(n1366), .IN3(n1361), .IN4(n1362), .IN5(
        n1377), .Q(n1353) );
  OA21X1 U1339 ( .IN1(n1378), .IN2(n1245), .IN3(n1359), .Q(n1377) );
  OR2X1 U1340 ( .IN1(n1350), .IN2(n1351), .Q(n1359) );
  OAI222X1 U1341 ( .IN1(n1379), .IN2(n1380), .IN3(n1381), .IN4(n1382), .IN5(
        n1383), .IN6(n1384), .QN(n1245) );
  OA22X1 U1342 ( .IN1(n1385), .IN2(n1386), .IN3(n1387), .IN4(n1388), .Q(n1383)
         );
  INVX0 U1343 ( .INP(n1389), .ZN(n1387) );
  OA22X1 U1344 ( .IN1(n1390), .IN2(n1391), .IN3(n1392), .IN4(n1393), .Q(n1386)
         );
  OA22X1 U1345 ( .IN1(n1394), .IN2(n1395), .IN3(n1396), .IN4(n1397), .Q(n1391)
         );
  OA21X1 U1346 ( .IN1(n1398), .IN2(n1399), .IN3(n1400), .Q(n1395) );
  NAND3X0 U1347 ( .IN1(n1401), .IN2(n1402), .IN3(n1403), .QN(n1400) );
  INVX0 U1348 ( .INP(n1404), .ZN(n1394) );
  AND2X1 U1349 ( .IN1(n1380), .IN2(n1379), .Q(n1381) );
  AO22X1 U1350 ( .IN1(n1405), .IN2(n1406), .IN3(n1407), .IN4(n1408), .Q(n1380)
         );
  NAND2X0 U1351 ( .IN1(n1409), .IN2(n1410), .QN(n1408) );
  INVX0 U1352 ( .INP(n1409), .ZN(n1406) );
  OA22X1 U1353 ( .IN1(n1411), .IN2(n1412), .IN3(n1413), .IN4(n1414), .Q(n1409)
         );
  AND2X1 U1354 ( .IN1(n1412), .IN2(n1411), .Q(n1414) );
  NOR2X0 U1355 ( .IN1(n1415), .IN2(n1416), .QN(n1412) );
  NOR2X0 U1356 ( .IN1(n1252), .IN2(n1246), .QN(n1378) );
  NAND4X0 U1357 ( .IN1(n1404), .IN2(n1402), .IN3(n1417), .IN4(n1418), .QN(
        n1246) );
  NOR3X0 U1358 ( .IN1(n1390), .IN2(n1385), .IN3(n1419), .QN(n1418) );
  NOR2X0 U1359 ( .IN1(n1403), .IN2(n1401), .QN(n1419) );
  NOR2X0 U1360 ( .IN1(n1389), .IN2(n1420), .QN(n1385) );
  AND2X1 U1361 ( .IN1(n1392), .IN2(n1393), .Q(n1390) );
  INVX0 U1362 ( .INP(n1384), .ZN(n1417) );
  AO221X1 U1363 ( .IN1(n1405), .IN2(n1407), .IN3(n1379), .IN4(n1382), .IN5(
        n1421), .Q(n1384) );
  AO22X1 U1364 ( .IN1(n1422), .IN2(n1423), .IN3(n1416), .IN4(n1415), .Q(n1421)
         );
  INVX0 U1365 ( .INP(n1424), .ZN(n1415) );
  INVX0 U1366 ( .INP(n1411), .ZN(n1422) );
  NAND2X0 U1367 ( .IN1(n1398), .IN2(n1399), .QN(n1402) );
  INVX0 U1368 ( .INP(n1425), .ZN(n1398) );
  NAND2X0 U1369 ( .IN1(n1396), .IN2(n1397), .QN(n1404) );
  NOR2X0 U1370 ( .IN1(n1250), .IN2(n1426), .QN(n1252) );
  OA221X1 U1371 ( .IN1(n1427), .IN2(n1428), .IN3(n1429), .IN4(n1430), .IN5(
        n1431), .Q(n1426) );
  OA221X1 U1372 ( .IN1(n1432), .IN2(n1433), .IN3(n1434), .IN4(n1435), .IN5(
        n1251), .Q(n1431) );
  NAND4X0 U1373 ( .IN1(n1436), .IN2(n1437), .IN3(n1438), .IN4(n1439), .QN(
        n1251) );
  NAND2X0 U1374 ( .IN1(n1440), .IN2(n1441), .QN(n1439) );
  AO221X1 U1375 ( .IN1(n1442), .IN2(n1443), .IN3(n1444), .IN4(n1445), .IN5(
        n1446), .Q(n1438) );
  OR2X1 U1376 ( .IN1(n1445), .IN2(n1444), .Q(n1443) );
  AO21X1 U1377 ( .IN1(n1447), .IN2(n1448), .IN3(n1449), .Q(n1445) );
  OA22X1 U1378 ( .IN1(n1447), .IN2(n1448), .IN3(n1450), .IN4(n1451), .Q(n1449)
         );
  NAND4X0 U1379 ( .IN1(n1452), .IN2(N70), .IN3(n1453), .IN4(n1454), .QN(n1437)
         );
  NAND3X0 U1380 ( .IN1(n1452), .IN2(n1455), .IN3(N89), .QN(n1436) );
  OR3X1 U1381 ( .IN1(N18), .IN2(N70), .IN3(n1453), .Q(n1455) );
  AOI221X1 U1382 ( .IN1(n1447), .IN2(n1448), .IN3(n1450), .IN4(n1451), .IN5(
        n1456), .QN(n1452) );
  AO21X1 U1383 ( .IN1(n1442), .IN2(n1444), .IN3(n1446), .Q(n1456) );
  NOR2X0 U1384 ( .IN1(n1441), .IN2(n1440), .QN(n1446) );
  INVX0 U1385 ( .INP(n1457), .ZN(n1444) );
  INVX0 U1386 ( .INP(n1458), .ZN(n1451) );
  OA22X1 U1387 ( .IN1(n1434), .IN2(n1459), .IN3(n1435), .IN4(n1460), .Q(n1250)
         );
  AND2X1 U1388 ( .IN1(n1459), .IN2(n1434), .Q(n1460) );
  OA22X1 U1389 ( .IN1(n1432), .IN2(n1461), .IN3(n1433), .IN4(n1462), .Q(n1459)
         );
  AND2X1 U1390 ( .IN1(n1461), .IN2(n1432), .Q(n1462) );
  OA22X1 U1391 ( .IN1(n1429), .IN2(n1463), .IN3(n1430), .IN4(n1464), .Q(n1461)
         );
  AND2X1 U1392 ( .IN1(n1463), .IN2(n1429), .Q(n1464) );
  AND2X1 U1393 ( .IN1(n1428), .IN2(n1427), .Q(n1463) );
  OA221X1 U1394 ( .IN1(n1355), .IN2(n1358), .IN3(n1373), .IN4(n1372), .IN5(
        n1465), .Q(n1352) );
  OA22X1 U1395 ( .IN1(n1376), .IN2(n1375), .IN3(n1368), .IN4(n1370), .Q(n1465)
         );
  OA222X1 U1396 ( .IN1(n1334), .IN2(n1335), .IN3(n1328), .IN4(n1466), .IN5(
        n1333), .IN6(n1467), .Q(n1313) );
  NAND4X0 U1397 ( .IN1(n1468), .IN2(n1469), .IN3(n1470), .IN4(n1471), .QN(
        N10576) );
  XOR3X1 U1398 ( .IN1(n1472), .IN2(n1473), .IN3(n1474), .Q(n1471) );
  AO21X1 U1399 ( .IN1(N164), .IN2(n1335), .IN3(n1475), .Q(n1474) );
  AO21X1 U1400 ( .IN1(N165), .IN2(n1335), .IN3(n1475), .Q(n1473) );
  AO221X1 U1401 ( .IN1(n1476), .IN2(n1477), .IN3(n1478), .IN4(n1479), .IN5(
        n1480), .Q(n1472) );
  MUX21X1 U1402 ( .IN1(n1481), .IN2(n1482), .S(n1483), .Q(n1480) );
  NOR2X0 U1403 ( .IN1(n1478), .IN2(n1484), .QN(n1482) );
  NOR2X0 U1404 ( .IN1(n1478), .IN2(n1485), .QN(n1481) );
  XOR2X1 U1405 ( .IN1(n1484), .IN2(keyinput18), .Q(n1485) );
  MUX21X1 U1406 ( .IN1(n1486), .IN2(n1487), .S(n1483), .Q(n1479) );
  NOR2X0 U1407 ( .IN1(n1486), .IN2(n1477), .QN(n1487) );
  INVX0 U1408 ( .INP(keyinput20), .ZN(n1477) );
  NAND3X0 U1409 ( .IN1(n1484), .IN2(n1478), .IN3(n1483), .QN(n1476) );
  NOR2X0 U1410 ( .IN1(N170), .IN2(n1488), .QN(n1483) );
  XOR2X1 U1411 ( .IN1(n1328), .IN2(n1333), .Q(n1478) );
  OA21X1 U1412 ( .IN1(N169), .IN2(n1475), .IN3(n1335), .Q(n1333) );
  OA21X1 U1413 ( .IN1(N168), .IN2(n1475), .IN3(n1335), .Q(n1328) );
  INVX0 U1414 ( .INP(n1486), .ZN(n1484) );
  XOR2X1 U1415 ( .IN1(n1316), .IN2(n1318), .Q(n1486) );
  OA21X1 U1416 ( .IN1(N167), .IN2(n1475), .IN3(n1335), .Q(n1318) );
  OA21X1 U1417 ( .IN1(N166), .IN2(n1475), .IN3(n1335), .Q(n1316) );
  XOR3X1 U1418 ( .IN1(n1489), .IN2(n1490), .IN3(n1491), .Q(n1470) );
  XNOR2X1 U1419 ( .IN1(n1355), .IN2(n1492), .Q(n1491) );
  NOR2X0 U1420 ( .IN1(keyinput15), .IN2(n1493), .QN(n1492) );
  XOR3X1 U1421 ( .IN1(n1368), .IN2(n1494), .IN3(n1361), .Q(n1493) );
  OA21X1 U1422 ( .IN1(N177), .IN2(n1475), .IN3(n1335), .Q(n1361) );
  XNOR2X1 U1423 ( .IN1(n1364), .IN2(n1373), .Q(n1494) );
  MUX21X1 U1424 ( .IN1(N138), .IN2(N180), .S(N18), .Q(n1373) );
  MUX21X1 U1425 ( .IN1(N135), .IN2(N178), .S(N18), .Q(n1364) );
  MUX21X1 U1426 ( .IN1(N144), .IN2(N179), .S(N18), .Q(n1368) );
  OA21X1 U1427 ( .IN1(N176), .IN2(n1475), .IN3(n1335), .Q(n1355) );
  MUX21X1 U1428 ( .IN1(n1495), .IN2(n1496), .S(N18), .Q(n1490) );
  XNOR2X1 U1429 ( .IN1(n1376), .IN2(N181), .Q(n1496) );
  XNOR2X1 U1430 ( .IN1(N141), .IN2(n1376), .Q(n1495) );
  MUX21X1 U1431 ( .IN1(N147), .IN2(N171), .S(N18), .Q(n1376) );
  XOR3X1 U1432 ( .IN1(n1340), .IN2(n1345), .IN3(n1351), .Q(n1489) );
  OA21X1 U1433 ( .IN1(N175), .IN2(n1475), .IN3(n1335), .Q(n1351) );
  INVX0 U1434 ( .INP(n1348), .ZN(n1345) );
  AO21X1 U1435 ( .IN1(N174), .IN2(n1335), .IN3(n1475), .Q(n1348) );
  INVX0 U1436 ( .INP(n1337), .ZN(n1340) );
  AO21X1 U1437 ( .IN1(N173), .IN2(n1335), .IN3(n1475), .Q(n1337) );
  XOR3X1 U1438 ( .IN1(n1497), .IN2(n1379), .IN3(n1498), .Q(n1469) );
  XOR3X1 U1439 ( .IN1(n1396), .IN2(n1499), .IN3(n1500), .Q(n1498) );
  MUX21X1 U1440 ( .IN1(n1501), .IN2(n1502), .S(N18), .Q(n1500) );
  XOR2X1 U1441 ( .IN1(N197), .IN2(n1403), .Q(n1502) );
  XOR2X1 U1442 ( .IN1(N115), .IN2(n1403), .Q(n1501) );
  MUX21X1 U1443 ( .IN1(N187), .IN2(N118), .S(n1454), .Q(n1403) );
  XOR2X1 U1444 ( .IN1(n1393), .IN2(n1389), .Q(n1499) );
  MUX21X1 U1445 ( .IN1(N47), .IN2(N193), .S(N18), .Q(n1389) );
  INVX0 U1446 ( .INP(n1503), .ZN(n1393) );
  MUX21X1 U1447 ( .IN1(N121), .IN2(N194), .S(N18), .Q(n1503) );
  INVX0 U1448 ( .INP(n1504), .ZN(n1396) );
  MUX21X1 U1449 ( .IN1(N94), .IN2(N195), .S(N18), .Q(n1504) );
  INVX0 U1450 ( .INP(n1505), .ZN(n1379) );
  MUX21X1 U1451 ( .IN1(N66), .IN2(N189), .S(N18), .Q(n1505) );
  XOR3X1 U1452 ( .IN1(n1424), .IN2(n1425), .IN3(n1506), .Q(n1497) );
  XOR2X1 U1453 ( .IN1(n1411), .IN2(n1405), .Q(n1506) );
  INVX0 U1454 ( .INP(n1410), .ZN(n1405) );
  MUX21X1 U1455 ( .IN1(N50), .IN2(N190), .S(N18), .Q(n1410) );
  MUX21X1 U1456 ( .IN1(N32), .IN2(N191), .S(N18), .Q(n1411) );
  MUX21X1 U1457 ( .IN1(N97), .IN2(N196), .S(N18), .Q(n1425) );
  MUX21X1 U1458 ( .IN1(N35), .IN2(N192), .S(N18), .Q(n1424) );
  XOR3X1 U1459 ( .IN1(n1458), .IN2(n1447), .IN3(n1507), .Q(n1468) );
  XOR2X1 U1460 ( .IN1(n1508), .IN2(n1509), .Q(n1507) );
  XOR3X1 U1461 ( .IN1(keyinput16), .IN2(n1441), .IN3(n1510), .Q(n1509) );
  XOR2X1 U1462 ( .IN1(n1432), .IN2(n1457), .Q(n1510) );
  MUX21X1 U1463 ( .IN1(N23), .IN2(N205), .S(N18), .Q(n1457) );
  MUX21X1 U1464 ( .IN1(N124), .IN2(N201), .S(N18), .Q(n1432) );
  MUX21X1 U1465 ( .IN1(N103), .IN2(N204), .S(N18), .Q(n1441) );
  XOR3X1 U1466 ( .IN1(n1428), .IN2(n1511), .IN3(n1512), .Q(n1508) );
  MUX21X1 U1467 ( .IN1(n1513), .IN2(n1514), .S(N18), .Q(n1512) );
  XNOR2X1 U1468 ( .IN1(N208), .IN2(n1453), .Q(n1514) );
  XNOR2X1 U1469 ( .IN1(N44), .IN2(n1453), .Q(n1513) );
  MUX21X1 U1470 ( .IN1(N41), .IN2(N198), .S(N18), .Q(n1453) );
  XOR2X1 U1471 ( .IN1(n1429), .IN2(n1434), .Q(n1511) );
  MUX21X1 U1472 ( .IN1(N100), .IN2(N200), .S(N18), .Q(n1434) );
  MUX21X1 U1473 ( .IN1(N127), .IN2(N202), .S(N18), .Q(n1429) );
  MUX21X1 U1474 ( .IN1(N130), .IN2(N203), .S(N18), .Q(n1428) );
  INVX0 U1475 ( .INP(n1515), .ZN(n1447) );
  MUX21X1 U1476 ( .IN1(N26), .IN2(N206), .S(N18), .Q(n1515) );
  MUX21X1 U1477 ( .IN1(N29), .IN2(N207), .S(N18), .Q(n1458) );
  NAND4X0 U1478 ( .IN1(n1516), .IN2(n1517), .IN3(n1518), .IN4(n1519), .QN(
        N10575) );
  XOR2X1 U1479 ( .IN1(n1520), .IN2(n1521), .Q(n1519) );
  XOR3X1 U1480 ( .IN1(n1315), .IN2(n1522), .IN3(n1321), .Q(n1521) );
  MUX21X1 U1481 ( .IN1(N112), .IN2(n1523), .S(N18), .Q(n1321) );
  INVX0 U1482 ( .INP(N257), .ZN(n1523) );
  MUX21X1 U1483 ( .IN1(n1524), .IN2(N267), .S(N18), .Q(n1522) );
  INVX0 U1484 ( .INP(N271), .ZN(n1524) );
  MUX21X1 U1485 ( .IN1(N88), .IN2(n1236), .S(N18), .Q(n1315) );
  INVX0 U1486 ( .INP(N260), .ZN(n1236) );
  XOR3X1 U1487 ( .IN1(n1331), .IN2(n1525), .IN3(n1526), .Q(n1520) );
  XOR2X1 U1488 ( .IN1(n1527), .IN2(n1326), .Q(n1526) );
  INVX0 U1489 ( .INP(n1466), .ZN(n1326) );
  MUX21X1 U1490 ( .IN1(N87), .IN2(n1528), .S(N18), .Q(n1466) );
  INVX0 U1491 ( .INP(N106), .ZN(n1528) );
  OA21X1 U1492 ( .IN1(n1334), .IN2(n1529), .IN3(n1530), .Q(n1527) );
  XOR2X1 U1493 ( .IN1(n1531), .IN2(keyinput6), .Q(n1530) );
  NAND2X0 U1494 ( .IN1(n1529), .IN2(n1334), .QN(n1531) );
  MUX21X1 U1495 ( .IN1(n1532), .IN2(N248), .S(N18), .Q(n1529) );
  INVX0 U1496 ( .INP(N114), .ZN(n1532) );
  MUX21X1 U1497 ( .IN1(N113), .IN2(n1253), .S(N18), .Q(n1334) );
  INVX0 U1498 ( .INP(N251), .ZN(n1253) );
  MUX21X1 U1499 ( .IN1(N245), .IN2(n1241), .S(N18), .Q(n1525) );
  INVX0 U1500 ( .INP(N263), .ZN(n1241) );
  INVX0 U1501 ( .INP(n1467), .ZN(n1331) );
  MUX21X1 U1502 ( .IN1(N111), .IN2(n1533), .S(N18), .Q(n1467) );
  INVX0 U1503 ( .INP(N254), .ZN(n1533) );
  XOR3X1 U1504 ( .IN1(n1382), .IN2(n1534), .IN3(n1535), .Q(n1518) );
  XOR3X1 U1505 ( .IN1(n1423), .IN2(n1536), .IN3(n1537), .Q(n1535) );
  MUX21X1 U1506 ( .IN1(n1538), .IN2(n1539), .S(N18), .Q(n1537) );
  XOR2X1 U1507 ( .IN1(n1540), .IN2(N337), .Q(n1539) );
  XOR2X1 U1508 ( .IN1(N58), .IN2(n1401), .Q(n1538) );
  INVX0 U1509 ( .INP(n1540), .ZN(n1401) );
  MUX21X1 U1510 ( .IN1(n1541), .IN2(N340), .S(N18), .Q(n1540) );
  INVX0 U1511 ( .INP(N77), .ZN(n1541) );
  XNOR2X1 U1512 ( .IN1(n1416), .IN2(n1407), .Q(n1536) );
  MUX21X1 U1513 ( .IN1(N361), .IN2(n1542), .S(n1454), .Q(n1407) );
  INVX0 U1514 ( .INP(N61), .ZN(n1542) );
  MUX21X1 U1515 ( .IN1(n1543), .IN2(N355), .S(N18), .Q(n1416) );
  INVX0 U1516 ( .INP(N79), .ZN(n1543) );
  INVX0 U1517 ( .INP(n1413), .ZN(n1423) );
  MUX21X1 U1518 ( .IN1(N60), .IN2(n1282), .S(N18), .Q(n1413) );
  INVX0 U1519 ( .INP(N358), .ZN(n1282) );
  XOR3X1 U1520 ( .IN1(n1388), .IN2(n1397), .IN3(n1544), .Q(n1534) );
  XOR2X1 U1521 ( .IN1(n1392), .IN2(n1545), .Q(n1544) );
  NOR2X0 U1522 ( .IN1(keyinput11), .IN2(n1399), .QN(n1545) );
  MUX21X1 U1523 ( .IN1(N343), .IN2(n1546), .S(n1454), .Q(n1399) );
  INVX0 U1524 ( .INP(N78), .ZN(n1546) );
  MUX21X1 U1525 ( .IN1(n1547), .IN2(N349), .S(N18), .Q(n1392) );
  INVX0 U1526 ( .INP(N81), .ZN(n1547) );
  MUX21X1 U1527 ( .IN1(N346), .IN2(n1548), .S(n1454), .Q(n1397) );
  INVX0 U1528 ( .INP(N59), .ZN(n1548) );
  INVX0 U1529 ( .INP(n1420), .ZN(n1388) );
  MUX21X1 U1530 ( .IN1(N80), .IN2(n1302), .S(N18), .Q(n1420) );
  INVX0 U1531 ( .INP(N352), .ZN(n1302) );
  MUX21X1 U1532 ( .IN1(N364), .IN2(n1549), .S(n1454), .Q(n1382) );
  INVX0 U1533 ( .INP(N62), .ZN(n1549) );
  XNOR3X1 U1534 ( .IN1(n1550), .IN2(n1551), .IN3(n1435), .Q(n1517) );
  MUX21X1 U1535 ( .IN1(N56), .IN2(n1552), .S(N18), .Q(n1435) );
  XOR3X1 U1536 ( .IN1(n1433), .IN2(n1427), .IN3(n1553), .Q(n1551) );
  XOR2X1 U1537 ( .IN1(n1430), .IN2(n1448), .Q(n1553) );
  INVX0 U1538 ( .INP(n1554), .ZN(n1448) );
  MUX21X1 U1539 ( .IN1(N76), .IN2(n1555), .S(N18), .Q(n1554) );
  MUX21X1 U1540 ( .IN1(N54), .IN2(n1556), .S(N18), .Q(n1430) );
  INVX0 U1541 ( .INP(N328), .ZN(n1556) );
  MUX21X1 U1542 ( .IN1(n1557), .IN2(N53), .S(n1454), .Q(n1427) );
  MUX21X1 U1543 ( .IN1(N55), .IN2(n1230), .S(N18), .Q(n1433) );
  XOR3X1 U1544 ( .IN1(n1440), .IN2(n1450), .IN3(n1558), .Q(n1550) );
  XNOR2X1 U1545 ( .IN1(n1559), .IN2(n1442), .Q(n1558) );
  MUX21X1 U1546 ( .IN1(n1560), .IN2(N319), .S(N18), .Q(n1442) );
  INVX0 U1547 ( .INP(N75), .ZN(n1560) );
  OA21X1 U1548 ( .IN1(n1561), .IN2(n1562), .IN3(n1563), .Q(n1559) );
  XOR2X1 U1549 ( .IN1(n1564), .IN2(keyinput9), .Q(n1563) );
  NAND2X0 U1550 ( .IN1(n1562), .IN2(n1561), .QN(n1564) );
  MUX21X1 U1551 ( .IN1(N70), .IN2(n1565), .S(N18), .Q(n1562) );
  MUX21X1 U1552 ( .IN1(n1566), .IN2(N307), .S(N18), .Q(n1561) );
  INVX0 U1553 ( .INP(N69), .ZN(n1566) );
  INVX0 U1554 ( .INP(n1567), .ZN(n1450) );
  MUX21X1 U1555 ( .IN1(N74), .IN2(n1568), .S(N18), .Q(n1567) );
  MUX21X1 U1556 ( .IN1(N73), .IN2(n1569), .S(N18), .Q(n1440) );
  XOR3X1 U1557 ( .IN1(n1342), .IN2(n1346), .IN3(n1570), .Q(n1516) );
  XNOR3X1 U1558 ( .IN1(n1571), .IN2(n1350), .IN3(n1572), .Q(n1570) );
  XOR3X1 U1559 ( .IN1(keyinput5), .IN2(n1573), .IN3(n1574), .Q(n1572) );
  XNOR2X1 U1560 ( .IN1(n1366), .IN2(n1370), .Q(n1574) );
  AO22X1 U1561 ( .IN1(N84), .IN2(n1575), .IN3(N18), .IN4(n1266), .Q(n1370) );
  INVX0 U1562 ( .INP(N283), .ZN(n1266) );
  AO22X1 U1563 ( .IN1(N85), .IN2(n1575), .IN3(N18), .IN4(n1576), .Q(n1366) );
  INVX0 U1564 ( .INP(N286), .ZN(n1576) );
  OA21X1 U1565 ( .IN1(N274), .IN2(n1454), .IN3(n1577), .Q(n1573) );
  NAND2X0 U1566 ( .IN1(N82), .IN2(n1575), .QN(n1577) );
  MUX21X1 U1567 ( .IN1(N86), .IN2(n1273), .S(N18), .Q(n1350) );
  INVX0 U1568 ( .INP(N296), .ZN(n1273) );
  XNOR3X1 U1569 ( .IN1(n1358), .IN2(n1362), .IN3(n1578), .Q(n1571) );
  XNOR2X1 U1570 ( .IN1(n1375), .IN2(n1372), .Q(n1578) );
  AO22X1 U1571 ( .IN1(N18), .IN2(n1579), .IN3(N83), .IN4(n1575), .Q(n1372) );
  INVX0 U1572 ( .INP(N280), .ZN(n1579) );
  AO21X1 U1573 ( .IN1(N65), .IN2(n1575), .IN3(n1580), .Q(n1375) );
  XOR2X1 U1574 ( .IN1(n1581), .IN2(keyinput2), .Q(n1580) );
  NAND2X0 U1575 ( .IN1(N18), .IN2(n1277), .QN(n1581) );
  INVX0 U1576 ( .INP(N277), .ZN(n1277) );
  XOR2X1 U1577 ( .IN1(N18), .IN2(keyinput1), .Q(n1575) );
  MUX21X1 U1578 ( .IN1(N64), .IN2(n1259), .S(N18), .Q(n1362) );
  INVX0 U1579 ( .INP(N289), .ZN(n1259) );
  MUX21X1 U1580 ( .IN1(N63), .IN2(n1582), .S(N18), .Q(n1358) );
  INVX0 U1581 ( .INP(N293), .ZN(n1582) );
  MUX21X1 U1582 ( .IN1(n1583), .IN2(N299), .S(N18), .Q(n1346) );
  INVX0 U1583 ( .INP(N109), .ZN(n1583) );
  MUX21X1 U1584 ( .IN1(n1584), .IN2(N303), .S(N18), .Q(n1342) );
  INVX0 U1585 ( .INP(N110), .ZN(n1584) );
  NAND4X0 U1586 ( .IN1(n1585), .IN2(n1586), .IN3(n1587), .IN4(n1588), .QN(
        N10574) );
  XOR3X1 U1587 ( .IN1(n1589), .IN2(n1590), .IN3(n1591), .Q(n1588) );
  XNOR3X1 U1588 ( .IN1(n1235), .IN2(n1239), .IN3(n1592), .Q(n1591) );
  XNOR2X1 U1589 ( .IN1(n1240), .IN2(n1238), .Q(n1592) );
  AOI21X1 U1590 ( .IN1(N216), .IN2(n1593), .IN3(n1594), .QN(n1238) );
  AOI21X1 U1591 ( .IN1(N214), .IN2(n1593), .IN3(n1594), .QN(n1240) );
  AOI21X1 U1592 ( .IN1(N215), .IN2(n1593), .IN3(n1594), .QN(n1239) );
  AO21X1 U1593 ( .IN1(N213), .IN2(n1335), .IN3(n1475), .Q(n1235) );
  AO21X1 U1594 ( .IN1(N211), .IN2(n1335), .IN3(n1475), .Q(n1590) );
  XOR2X1 U1595 ( .IN1(n1595), .IN2(n1596), .Q(n1589) );
  NOR2X0 U1596 ( .IN1(n1488), .IN2(n1254), .QN(n1596) );
  AO21X1 U1597 ( .IN1(N209), .IN2(n1593), .IN3(n1594), .Q(n1254) );
  MUX21X1 U1598 ( .IN1(n1593), .IN2(n1475), .S(keyinput0), .Q(n1594) );
  INVX0 U1599 ( .INP(n1488), .ZN(n1593) );
  NAND2X0 U1600 ( .IN1(N18), .IN2(n1335), .QN(n1488) );
  AO21X1 U1601 ( .IN1(N212), .IN2(n1335), .IN3(n1475), .Q(n1595) );
  XOR3X1 U1602 ( .IN1(n1597), .IN2(n1598), .IN3(n1599), .Q(n1587) );
  XNOR2X1 U1603 ( .IN1(n1267), .IN2(n1600), .Q(n1599) );
  OA21X1 U1604 ( .IN1(n1601), .IN2(n1265), .IN3(n1602), .Q(n1600) );
  XOR2X1 U1605 ( .IN1(n1603), .IN2(keyinput7), .Q(n1602) );
  NAND2X0 U1606 ( .IN1(n1601), .IN2(n1265), .QN(n1603) );
  MUX21X1 U1607 ( .IN1(N135), .IN2(N158), .S(N18), .Q(n1265) );
  INVX0 U1608 ( .INP(n1258), .ZN(n1601) );
  AO21X1 U1609 ( .IN1(N157), .IN2(n1335), .IN3(n1475), .Q(n1258) );
  MUX21X1 U1610 ( .IN1(N144), .IN2(N159), .S(N18), .Q(n1267) );
  XOR3X1 U1611 ( .IN1(n1275), .IN2(n1270), .IN3(n1604), .Q(n1598) );
  XOR2X1 U1612 ( .IN1(n1272), .IN2(n1274), .Q(n1604) );
  OA21X1 U1613 ( .IN1(N156), .IN2(n1475), .IN3(n1335), .Q(n1274) );
  OA21X1 U1614 ( .IN1(N155), .IN2(n1475), .IN3(n1335), .Q(n1272) );
  AOI21X1 U1615 ( .IN1(N153), .IN2(n1335), .IN3(n1475), .QN(n1270) );
  AOI21X1 U1616 ( .IN1(N154), .IN2(n1335), .IN3(n1475), .QN(n1275) );
  AND2X1 U1617 ( .IN1(n1335), .IN2(n1454), .Q(n1475) );
  NAND2X0 U1618 ( .IN1(N9), .IN2(N12), .QN(n1335) );
  XOR2X1 U1619 ( .IN1(n1269), .IN2(n1605), .Q(n1597) );
  MUX21X1 U1620 ( .IN1(n1606), .IN2(n1607), .S(N18), .Q(n1605) );
  XOR2X1 U1621 ( .IN1(n1276), .IN2(N161), .Q(n1607) );
  XOR2X1 U1622 ( .IN1(n1276), .IN2(N141), .Q(n1606) );
  MUX21X1 U1623 ( .IN1(N147), .IN2(N151), .S(N18), .Q(n1276) );
  MUX21X1 U1624 ( .IN1(N138), .IN2(N160), .S(N18), .Q(n1269) );
  XOR3X1 U1625 ( .IN1(n1306), .IN2(n1304), .IN3(n1608), .Q(n1586) );
  XOR3X1 U1626 ( .IN1(n1281), .IN2(n1309), .IN3(n1609), .Q(n1608) );
  NAND2X0 U1627 ( .IN1(n1610), .IN2(n1611), .QN(n1609) );
  XOR2X1 U1628 ( .IN1(n1612), .IN2(keyinput21), .Q(n1611) );
  NAND3X0 U1629 ( .IN1(n1613), .IN2(n1614), .IN3(n1615), .QN(n1612) );
  MUX21X1 U1630 ( .IN1(n1616), .IN2(n1617), .S(n1614), .Q(n1610) );
  INVX0 U1631 ( .INP(n1618), .ZN(n1614) );
  MUX21X1 U1632 ( .IN1(n1619), .IN2(n1620), .S(N18), .Q(n1618) );
  XOR2X1 U1633 ( .IN1(n1299), .IN2(N227), .Q(n1620) );
  XOR2X1 U1634 ( .IN1(n1299), .IN2(N115), .Q(n1619) );
  MUX21X1 U1635 ( .IN1(N118), .IN2(N217), .S(N18), .Q(n1299) );
  OR2X1 U1636 ( .IN1(n1615), .IN2(n1613), .Q(n1617) );
  XNOR2X1 U1637 ( .IN1(n1613), .IN2(n1615), .Q(n1616) );
  XNOR2X1 U1638 ( .IN1(n1301), .IN2(n1234), .Q(n1615) );
  INVX0 U1639 ( .INP(n1293), .ZN(n1234) );
  MUX21X1 U1640 ( .IN1(N224), .IN2(N121), .S(n1454), .Q(n1293) );
  MUX21X1 U1641 ( .IN1(N47), .IN2(N223), .S(N18), .Q(n1301) );
  XOR2X1 U1642 ( .IN1(n1298), .IN2(n1300), .Q(n1613) );
  INVX0 U1643 ( .INP(n1621), .ZN(n1300) );
  MUX21X1 U1644 ( .IN1(N94), .IN2(N225), .S(N18), .Q(n1621) );
  MUX21X1 U1645 ( .IN1(N97), .IN2(N226), .S(N18), .Q(n1298) );
  MUX21X1 U1646 ( .IN1(N35), .IN2(N222), .S(N18), .Q(n1309) );
  MUX21X1 U1647 ( .IN1(N32), .IN2(N221), .S(N18), .Q(n1281) );
  MUX21X1 U1648 ( .IN1(N66), .IN2(N219), .S(N18), .Q(n1304) );
  MUX21X1 U1649 ( .IN1(N50), .IN2(N220), .S(N18), .Q(n1306) );
  XOR3X1 U1650 ( .IN1(n1622), .IN2(n1623), .IN3(n1624), .Q(n1585) );
  XOR3X1 U1651 ( .IN1(n1231), .IN2(n1625), .IN3(n1626), .Q(n1624) );
  NAND2X0 U1652 ( .IN1(n1627), .IN2(keyinput25), .QN(n1626) );
  XOR2X1 U1653 ( .IN1(n1628), .IN2(n1629), .Q(n1627) );
  XNOR3X1 U1654 ( .IN1(n1630), .IN2(n1631), .IN3(n1632), .Q(n1629) );
  MUX21X1 U1655 ( .IN1(n1633), .IN2(n1634), .S(N18), .Q(n1632) );
  XOR2X1 U1656 ( .IN1(n1635), .IN2(N239), .Q(n1634) );
  XOR2X1 U1657 ( .IN1(n1635), .IN2(N44), .Q(n1633) );
  XOR3X1 U1658 ( .IN1(keyinput14), .IN2(n1636), .IN3(n1637), .Q(n1628) );
  XOR2X1 U1659 ( .IN1(n965), .IN2(n1638), .Q(N10353) );
  XOR2X1 U1660 ( .IN1(n966), .IN2(n1639), .Q(N10352) );
  OA21X1 U1661 ( .IN1(n1640), .IN2(n1638), .IN3(n963), .Q(n1639) );
  XOR2X1 U1662 ( .IN1(n1290), .IN2(n1641), .Q(N10351) );
  OA21X1 U1663 ( .IN1(n972), .IN2(n1638), .IN3(n1229), .Q(n1641) );
  MUX21X1 U1664 ( .IN1(n1642), .IN2(n1643), .S(n1638), .Q(N10350) );
  INVX0 U1665 ( .INP(n1228), .ZN(n1638) );
  AO21X1 U1666 ( .IN1(N367), .IN2(n956), .IN3(n955), .Q(n1228) );
  AO22X1 U1667 ( .IN1(n1636), .IN2(n1569), .IN3(n923), .IN4(n1644), .Q(n955)
         );
  NAND3X0 U1668 ( .IN1(n1645), .IN2(n1646), .IN3(n1647), .QN(n1644) );
  NAND2X0 U1669 ( .IN1(n1648), .IN2(n938), .QN(n1647) );
  AND2X1 U1670 ( .IN1(n940), .IN2(n923), .Q(n956) );
  NOR2X0 U1671 ( .IN1(n939), .IN2(n927), .QN(n940) );
  INVX0 U1672 ( .INP(n1648), .ZN(n927) );
  NOR2X0 U1673 ( .IN1(n1291), .IN2(n1649), .QN(n1643) );
  NOR3X0 U1674 ( .IN1(n1650), .IN2(n962), .IN3(n1651), .QN(n1649) );
  OA21X1 U1675 ( .IN1(n1650), .IN2(n1651), .IN3(n962), .Q(n1291) );
  NOR2X0 U1676 ( .IN1(n1229), .IN2(n1290), .QN(n1650) );
  XNOR2X1 U1677 ( .IN1(n962), .IN2(n1652), .Q(n1642) );
  OA21X1 U1678 ( .IN1(n972), .IN2(n1290), .IN3(n973), .Q(n1652) );
  AO22X1 U1679 ( .IN1(n1651), .IN2(keyinput10), .IN3(n1653), .IN4(n1654), .Q(
        n1290) );
  NAND2X0 U1680 ( .IN1(keyinput10), .IN2(n1230), .QN(n1654) );
  INVX0 U1681 ( .INP(n1231), .ZN(n1653) );
  INVX0 U1682 ( .INP(n973), .ZN(n1651) );
  NAND2X0 U1683 ( .IN1(n1231), .IN2(n1230), .QN(n973) );
  INVX0 U1684 ( .INP(N331), .ZN(n1230) );
  MUX21X1 U1685 ( .IN1(N124), .IN2(N232), .S(N18), .Q(n1231) );
  NOR2X0 U1686 ( .IN1(n961), .IN2(n967), .QN(n972) );
  NOR2X0 U1687 ( .IN1(n965), .IN2(n966), .QN(n967) );
  NAND2X0 U1688 ( .IN1(n976), .IN2(n963), .QN(n965) );
  INVX0 U1689 ( .INP(n1640), .ZN(n976) );
  NOR2X0 U1690 ( .IN1(n1557), .IN2(n1622), .QN(n1640) );
  INVX0 U1691 ( .INP(n1229), .ZN(n961) );
  OA22X1 U1692 ( .IN1(n1623), .IN2(N328), .IN3(n963), .IN4(n966), .Q(n1229) );
  XNOR2X1 U1693 ( .IN1(n1623), .IN2(N328), .Q(n966) );
  NAND2X0 U1694 ( .IN1(n1622), .IN2(n1557), .QN(n963) );
  INVX0 U1695 ( .INP(N325), .ZN(n1557) );
  MUX21X1 U1696 ( .IN1(N130), .IN2(N234), .S(N18), .Q(n1622) );
  INVX0 U1697 ( .INP(n1655), .ZN(n1623) );
  MUX21X1 U1698 ( .IN1(N127), .IN2(N233), .S(N18), .Q(n1655) );
  OA21X1 U1699 ( .IN1(n1552), .IN2(n1625), .IN3(n1226), .Q(n962) );
  NAND2X0 U1700 ( .IN1(n1625), .IN2(n1552), .QN(n1226) );
  MUX21X1 U1701 ( .IN1(N100), .IN2(N231), .S(N18), .Q(n1625) );
  INVX0 U1702 ( .INP(N334), .ZN(n1552) );
  XNOR2X1 U1703 ( .IN1(n932), .IN2(n1656), .Q(N10112) );
  OA21X1 U1704 ( .IN1(n1657), .IN2(n952), .IN3(n1658), .Q(n1656) );
  XOR2X1 U1705 ( .IN1(n947), .IN2(n1659), .Q(N10111) );
  NOR2X0 U1706 ( .IN1(n1660), .IN2(n938), .QN(n1659) );
  AO22X1 U1707 ( .IN1(n1631), .IN2(n1568), .IN3(n946), .IN4(n932), .Q(n938) );
  AO21X1 U1708 ( .IN1(n1661), .IN2(n930), .IN3(n1662), .Q(N10110) );
  XOR2X1 U1709 ( .IN1(n1663), .IN2(keyinput26), .Q(n1662) );
  OR2X1 U1710 ( .IN1(n1661), .IN2(n930), .Q(n1663) );
  AO21X1 U1711 ( .IN1(n1660), .IN2(n924), .IN3(n937), .Q(n1661) );
  NAND3X0 U1712 ( .IN1(n1664), .IN2(n1665), .IN3(n1666), .QN(n937) );
  NAND3X0 U1713 ( .IN1(n924), .IN2(n1568), .IN3(n1631), .QN(n1666) );
  XNOR2X1 U1714 ( .IN1(n1667), .IN2(n923), .Q(N10109) );
  XOR2X1 U1715 ( .IN1(n1569), .IN2(n1636), .Q(n923) );
  MUX21X1 U1716 ( .IN1(N103), .IN2(N235), .S(N18), .Q(n1636) );
  INVX0 U1717 ( .INP(N322), .ZN(n1569) );
  AOI21X1 U1718 ( .IN1(n1648), .IN2(n1660), .IN3(n941), .QN(n1667) );
  NAND4X0 U1719 ( .IN1(n1668), .IN2(n1669), .IN3(n1645), .IN4(n1646), .QN(n941) );
  INVX0 U1720 ( .INP(n1670), .ZN(n1646) );
  OR2X1 U1721 ( .IN1(n930), .IN2(n1665), .Q(n1645) );
  OR2X1 U1722 ( .IN1(n1664), .IN2(n930), .Q(n1669) );
  NAND3X0 U1723 ( .IN1(n932), .IN2(n924), .IN3(n946), .QN(n1664) );
  INVX0 U1724 ( .INP(n1658), .ZN(n946) );
  NAND3X0 U1725 ( .IN1(n1631), .IN2(n1568), .IN3(n1648), .QN(n1668) );
  INVX0 U1726 ( .INP(N313), .ZN(n1568) );
  NOR2X0 U1727 ( .IN1(n952), .IN2(n939), .QN(n1660) );
  NAND2X0 U1728 ( .IN1(n919), .IN2(n932), .QN(n939) );
  XNOR2X1 U1729 ( .IN1(n1631), .IN2(N313), .Q(n932) );
  MUX21X1 U1730 ( .IN1(N29), .IN2(N238), .S(N18), .Q(n1631) );
  INVX0 U1731 ( .INP(N367), .ZN(n952) );
  NOR2X0 U1732 ( .IN1(n947), .IN2(n930), .QN(n1648) );
  AO21X1 U1733 ( .IN1(N319), .IN2(n1637), .IN3(n1670), .Q(n930) );
  NOR2X0 U1734 ( .IN1(n1637), .IN2(N319), .QN(n1670) );
  INVX0 U1735 ( .INP(n1671), .ZN(n1637) );
  MUX21X1 U1736 ( .IN1(N23), .IN2(N236), .S(N18), .Q(n1671) );
  INVX0 U1737 ( .INP(n924), .ZN(n947) );
  OA21X1 U1738 ( .IN1(n1555), .IN2(n1630), .IN3(n1665), .Q(n924) );
  NAND2X0 U1739 ( .IN1(n1630), .IN2(n1555), .QN(n1665) );
  MUX21X1 U1740 ( .IN1(N26), .IN2(N237), .S(N18), .Q(n1630) );
  INVX0 U1741 ( .INP(N316), .ZN(n1555) );
  XOR2X1 U1742 ( .IN1(N367), .IN2(n919), .Q(N10025) );
  INVX0 U1743 ( .INP(n1657), .ZN(n919) );
  NAND2X0 U1744 ( .IN1(n934), .IN2(n1658), .QN(n1657) );
  NAND3X0 U1745 ( .IN1(n1672), .IN2(n1454), .IN3(n1635), .QN(n1658) );
  OR2X1 U1746 ( .IN1(n1672), .IN2(n1635), .Q(n934) );
  MUX21X1 U1747 ( .IN1(N41), .IN2(N229), .S(N18), .Q(n1635) );
  NAND2X0 U1748 ( .IN1(n1673), .IN2(n1454), .QN(n1672) );
  INVX0 U1749 ( .INP(N18), .ZN(n1454) );
  XOR2X1 U1750 ( .IN1(n1565), .IN2(keyinput4), .Q(n1673) );
  INVX0 U1751 ( .INP(N310), .ZN(n1565) );
endmodule

