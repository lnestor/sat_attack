
module c1908 ( N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, 
        N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, 
        N85, N88, N91, N94, N99, N104, N2753, N2754, N2755, N2756, N2762, 
        N2767, N2768, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, 
        N2787, N2811, N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43,
         N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88,
         N91, N94, N99, N104, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781,
         N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888,
         N2889, N2890, N2891, N2892, N2899;
  wire   n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766;

  NOR2X0 U411 ( .IN1(n402), .IN2(n403), .QN(N2899) );
  XOR3X1 U412 ( .IN1(N1), .IN2(n404), .IN3(n405), .Q(n403) );
  NAND2X0 U413 ( .IN1(keyinput15), .IN2(n406), .QN(n405) );
  NAND2X0 U414 ( .IN1(n407), .IN2(keyinput48), .QN(n404) );
  XOR3X1 U415 ( .IN1(keyinput120), .IN2(n408), .IN3(n409), .Q(n407) );
  NAND2X0 U416 ( .IN1(n410), .IN2(N79), .QN(n409) );
  OA21X1 U417 ( .IN1(n411), .IN2(n412), .IN3(keyinput123), .Q(n408) );
  XNOR2X1 U418 ( .IN1(keyinput68), .IN2(n413), .Q(n412) );
  XOR2X1 U419 ( .IN1(keyinput6), .IN2(n414), .Q(n402) );
  AO21X1 U420 ( .IN1(n415), .IN2(n416), .IN3(n417), .Q(N2892) );
  XNOR2X1 U421 ( .IN1(keyinput126), .IN2(n418), .Q(n417) );
  NOR2X0 U422 ( .IN1(n415), .IN2(n419), .QN(n418) );
  AOI21X1 U423 ( .IN1(N66), .IN2(N91), .IN3(n420), .QN(n419) );
  AO21X1 U424 ( .IN1(N104), .IN2(n421), .IN3(n422), .Q(n416) );
  AOI21X1 U425 ( .IN1(n423), .IN2(n424), .IN3(n425), .QN(n415) );
  XOR2X1 U426 ( .IN1(n426), .IN2(keyinput118), .Q(n425) );
  NAND3X0 U427 ( .IN1(n427), .IN2(n420), .IN3(n428), .QN(n426) );
  INVX0 U428 ( .INP(n423), .ZN(n427) );
  NAND2X0 U429 ( .IN1(n428), .IN2(n420), .QN(n424) );
  NOR2X0 U430 ( .IN1(n429), .IN2(n422), .QN(n423) );
  XOR2X1 U431 ( .IN1(keyinput72), .IN2(n430), .Q(n429) );
  OA21X1 U432 ( .IN1(n431), .IN2(n432), .IN3(n433), .Q(n430) );
  XOR2X1 U433 ( .IN1(n434), .IN2(keyinput67), .Q(n433) );
  NAND2X0 U434 ( .IN1(n432), .IN2(n431), .QN(n434) );
  XOR2X1 U435 ( .IN1(n435), .IN2(n436), .Q(n432) );
  XOR3X1 U436 ( .IN1(n437), .IN2(n438), .IN3(n439), .Q(n435) );
  XNOR2X1 U437 ( .IN1(n440), .IN2(n441), .Q(N2891) );
  NOR3X0 U438 ( .IN1(n442), .IN2(keyinput125), .IN3(n420), .QN(n441) );
  XOR2X1 U439 ( .IN1(keyinput3), .IN2(n443), .Q(n442) );
  NOR2X0 U440 ( .IN1(n444), .IN2(n445), .QN(n443) );
  OA21X1 U441 ( .IN1(n446), .IN2(n447), .IN3(n448), .Q(n440) );
  XOR2X1 U442 ( .IN1(n449), .IN2(keyinput117), .Q(n448) );
  NAND3X0 U443 ( .IN1(n450), .IN2(n420), .IN3(n447), .QN(n449) );
  AO21X1 U444 ( .IN1(N104), .IN2(n445), .IN3(n451), .Q(n447) );
  XOR2X1 U445 ( .IN1(n452), .IN2(n453), .Q(n451) );
  NAND2X0 U446 ( .IN1(n454), .IN2(keyinput50), .QN(n452) );
  XOR2X1 U447 ( .IN1(n455), .IN2(n456), .Q(n454) );
  NOR2X0 U448 ( .IN1(n457), .IN2(keyinput60), .QN(n456) );
  AND2X1 U449 ( .IN1(n420), .IN2(n450), .Q(n446) );
  NOR2X0 U450 ( .IN1(n414), .IN2(n458), .QN(N2890) );
  XOR2X1 U451 ( .IN1(n459), .IN2(n460), .Q(n458) );
  NAND2X0 U452 ( .IN1(n410), .IN2(n461), .QN(n459) );
  NOR2X0 U453 ( .IN1(n414), .IN2(n462), .QN(N2889) );
  OA21X1 U454 ( .IN1(n463), .IN2(n464), .IN3(n465), .Q(n462) );
  XOR2X1 U455 ( .IN1(keyinput121), .IN2(n466), .Q(n465) );
  AND2X1 U456 ( .IN1(n464), .IN2(n463), .Q(n466) );
  AND2X1 U457 ( .IN1(n410), .IN2(N85), .Q(n463) );
  NOR2X0 U458 ( .IN1(n414), .IN2(n467), .QN(N2888) );
  OA21X1 U459 ( .IN1(n468), .IN2(n469), .IN3(n470), .Q(n467) );
  XOR2X1 U460 ( .IN1(n471), .IN2(keyinput124), .Q(n470) );
  NAND2X0 U461 ( .IN1(n468), .IN2(n469), .QN(n471) );
  XOR2X1 U462 ( .IN1(n472), .IN2(keyinput119), .Q(n468) );
  NAND2X0 U463 ( .IN1(n410), .IN2(N82), .QN(n472) );
  NOR2X0 U464 ( .IN1(n414), .IN2(n473), .QN(N2887) );
  XOR3X1 U465 ( .IN1(keyinput127), .IN2(n474), .IN3(n475), .Q(n473) );
  NOR2X0 U466 ( .IN1(keyinput122), .IN2(n476), .QN(n475) );
  XOR3X1 U467 ( .IN1(n477), .IN2(n478), .IN3(n479), .Q(n476) );
  XNOR2X1 U468 ( .IN1(n480), .IN2(n481), .Q(n479) );
  NAND2X0 U469 ( .IN1(keyinput28), .IN2(n482), .QN(n478) );
  XOR3X1 U470 ( .IN1(keyinput83), .IN2(keyinput76), .IN3(N40), .Q(n477) );
  AND2X1 U471 ( .IN1(N76), .IN2(n410), .Q(n474) );
  NOR2X0 U472 ( .IN1(n483), .IN2(n484), .QN(N2886) );
  XOR3X1 U473 ( .IN1(n485), .IN2(n486), .IN3(n487), .Q(n484) );
  NAND2X0 U474 ( .IN1(n410), .IN2(n488), .QN(n486) );
  NOR2X0 U475 ( .IN1(n489), .IN2(n490), .QN(n410) );
  OA21X1 U476 ( .IN1(n491), .IN2(n492), .IN3(n493), .Q(n485) );
  XOR2X1 U477 ( .IN1(keyinput66), .IN2(n494), .Q(n493) );
  AND2X1 U478 ( .IN1(n491), .IN2(n492), .Q(n494) );
  XNOR2X1 U479 ( .IN1(n495), .IN2(n496), .Q(n492) );
  NAND2X0 U480 ( .IN1(keyinput59), .IN2(n497), .QN(n495) );
  XNOR2X1 U481 ( .IN1(n414), .IN2(keyinput5), .Q(n483) );
  NOR2X0 U482 ( .IN1(n420), .IN2(N99), .QN(n414) );
  AND2X1 U483 ( .IN1(n498), .IN2(n499), .Q(N2811) );
  NAND4X0 U484 ( .IN1(N99), .IN2(n500), .IN3(n490), .IN4(n501), .QN(n499) );
  NOR4X0 U485 ( .IN1(N104), .IN2(n502), .IN3(n503), .IN4(n504), .QN(n501) );
  NOR2X0 U486 ( .IN1(n505), .IN2(n506), .QN(n504) );
  INVX0 U487 ( .INP(n507), .ZN(n506) );
  OA22X1 U488 ( .IN1(n508), .IN2(n509), .IN3(n510), .IN4(n511), .Q(n505) );
  OA21X1 U489 ( .IN1(n512), .IN2(n513), .IN3(n514), .Q(n508) );
  NOR4X0 U490 ( .IN1(n515), .IN2(n511), .IN3(n509), .IN4(n516), .QN(n503) );
  OA22X1 U491 ( .IN1(n517), .IN2(n518), .IN3(n519), .IN4(n520), .Q(n515) );
  AOI21X1 U492 ( .IN1(n521), .IN2(n522), .IN3(n523), .QN(n519) );
  NOR2X0 U493 ( .IN1(n524), .IN2(n525), .QN(n517) );
  NOR2X0 U494 ( .IN1(n428), .IN2(n450), .QN(n490) );
  NAND4X0 U495 ( .IN1(n526), .IN2(n527), .IN3(n528), .IN4(n529), .QN(n450) );
  AND4X1 U496 ( .IN1(n530), .IN2(n531), .IN3(n532), .IN4(n533), .Q(n529) );
  AND2X1 U497 ( .IN1(n534), .IN2(n535), .Q(n528) );
  XNOR2X1 U498 ( .IN1(keyinput97), .IN2(n536), .Q(n527) );
  XOR2X1 U499 ( .IN1(n537), .IN2(keyinput94), .Q(n526) );
  NAND4X0 U500 ( .IN1(n538), .IN2(n539), .IN3(n540), .IN4(n541), .QN(n428) );
  NOR4X0 U501 ( .IN1(n542), .IN2(n543), .IN3(n544), .IN4(n545), .QN(n541) );
  XOR2X1 U502 ( .IN1(n546), .IN2(keyinput98), .Q(n545) );
  AND2X1 U503 ( .IN1(n547), .IN2(n548), .Q(n540) );
  XNOR2X1 U504 ( .IN1(n549), .IN2(keyinput99), .Q(n500) );
  NAND4X0 U505 ( .IN1(n550), .IN2(n507), .IN3(n551), .IN4(n552), .QN(n549) );
  NOR3X0 U506 ( .IN1(n518), .IN2(n520), .IN3(n516), .QN(n507) );
  INVX0 U507 ( .INP(n553), .ZN(n520) );
  INVX0 U508 ( .INP(n554), .ZN(n518) );
  XNOR2X1 U509 ( .IN1(n555), .IN2(keyinput93), .Q(n498) );
  OR3X1 U510 ( .IN1(N104), .IN2(N99), .IN3(n502), .Q(n555) );
  AND4X1 U511 ( .IN1(n556), .IN2(n557), .IN3(n558), .IN4(n559), .Q(n502) );
  NOR4X0 U512 ( .IN1(n560), .IN2(n561), .IN3(n562), .IN4(n563), .QN(n559) );
  MUX21X1 U513 ( .IN1(n564), .IN2(n565), .S(N76), .Q(n563) );
  AND2X1 U514 ( .IN1(n566), .IN2(keyinput10), .Q(n565) );
  MUX21X1 U515 ( .IN1(n567), .IN2(n568), .S(n566), .Q(n564) );
  NAND2X0 U516 ( .IN1(keyinput10), .IN2(n567), .QN(n568) );
  INVX0 U517 ( .INP(keyinput86), .ZN(n567) );
  XOR3X1 U518 ( .IN1(keyinput89), .IN2(n488), .IN3(n569), .Q(n562) );
  NOR2X0 U519 ( .IN1(n570), .IN2(keyinput35), .QN(n569) );
  XOR2X1 U520 ( .IN1(n571), .IN2(n572), .Q(n561) );
  NOR2X0 U521 ( .IN1(n573), .IN2(keyinput12), .QN(n571) );
  NOR3X0 U522 ( .IN1(n550), .IN2(n574), .IN3(n575), .QN(n558) );
  NAND2X0 U523 ( .IN1(n576), .IN2(n577), .QN(n557) );
  XOR2X1 U524 ( .IN1(keyinput11), .IN2(N82), .Q(n576) );
  XOR3X1 U525 ( .IN1(keyinput82), .IN2(n461), .IN3(n578), .Q(n556) );
  XNOR3X1 U526 ( .IN1(keyinput102), .IN2(N40), .IN3(n544), .Q(N2787) );
  AND3X1 U527 ( .IN1(n579), .IN2(n580), .IN3(n522), .Q(n544) );
  XNOR3X1 U528 ( .IN1(keyinput116), .IN2(N37), .IN3(n539), .Q(N2786) );
  NAND4X0 U529 ( .IN1(n553), .IN2(n580), .IN3(n521), .IN4(n560), .QN(n539) );
  XOR3X1 U530 ( .IN1(keyinput101), .IN2(N34), .IN3(n548), .Q(N2785) );
  NAND3X0 U531 ( .IN1(n525), .IN2(n523), .IN3(n580), .QN(n548) );
  AO21X1 U532 ( .IN1(n543), .IN2(n581), .IN3(n582), .Q(N2784) );
  XOR2X1 U533 ( .IN1(keyinput113), .IN2(n583), .Q(n582) );
  NOR2X0 U534 ( .IN1(n543), .IN2(n581), .QN(n583) );
  AND3X1 U535 ( .IN1(n523), .IN2(n580), .IN3(n524), .Q(n543) );
  NOR3X0 U536 ( .IN1(n510), .IN2(n584), .IN3(n511), .QN(n580) );
  INVX0 U537 ( .INP(n552), .ZN(n511) );
  NOR2X0 U538 ( .IN1(n512), .IN2(n575), .QN(n552) );
  XOR2X1 U539 ( .IN1(n585), .IN2(keyinput90), .Q(n512) );
  XOR2X1 U540 ( .IN1(n546), .IN2(n586), .Q(N2783) );
  NAND2X0 U541 ( .IN1(keyinput108), .IN2(N25), .QN(n586) );
  NAND4X0 U542 ( .IN1(n522), .IN2(n587), .IN3(n588), .IN4(n579), .QN(n546) );
  NOR2X0 U543 ( .IN1(n584), .IN2(n514), .QN(n588) );
  XNOR2X1 U544 ( .IN1(N22), .IN2(n536), .Q(N2782) );
  NAND4X0 U545 ( .IN1(n589), .IN2(n554), .IN3(n590), .IN4(n591), .QN(n536) );
  XOR2X1 U546 ( .IN1(n592), .IN2(n535), .Q(N2781) );
  NAND4X0 U547 ( .IN1(n589), .IN2(n553), .IN3(n521), .IN4(n560), .QN(n535) );
  NAND2X0 U548 ( .IN1(n593), .IN2(n594), .QN(N2780) );
  XOR2X1 U549 ( .IN1(keyinput107), .IN2(n595), .Q(n594) );
  NOR2X0 U550 ( .IN1(N16), .IN2(n596), .QN(n595) );
  XOR2X1 U551 ( .IN1(n534), .IN2(keyinput100), .Q(n596) );
  XOR2X1 U552 ( .IN1(keyinput112), .IN2(n597), .Q(n593) );
  NOR2X0 U553 ( .IN1(n598), .IN2(n599), .QN(n597) );
  XNOR2X1 U554 ( .IN1(keyinput100), .IN2(n534), .Q(n599) );
  NAND3X0 U555 ( .IN1(n525), .IN2(n523), .IN3(n589), .QN(n534) );
  INVX0 U556 ( .INP(N16), .ZN(n598) );
  XOR2X1 U557 ( .IN1(n600), .IN2(keyinput115), .Q(N2779) );
  NAND2X0 U558 ( .IN1(n601), .IN2(n602), .QN(n600) );
  XOR2X1 U559 ( .IN1(keyinput106), .IN2(n603), .Q(n602) );
  NOR2X0 U560 ( .IN1(N13), .IN2(n533), .QN(n603) );
  XOR2X1 U561 ( .IN1(n604), .IN2(keyinput111), .Q(n601) );
  NAND2X0 U562 ( .IN1(N13), .IN2(n533), .QN(n604) );
  NAND3X0 U563 ( .IN1(n523), .IN2(n524), .IN3(n589), .QN(n533) );
  AND2X1 U564 ( .IN1(n605), .IN2(n587), .Q(n589) );
  INVX0 U565 ( .INP(n509), .ZN(n587) );
  NAND2X0 U566 ( .IN1(n551), .IN2(n606), .QN(n509) );
  INVX0 U567 ( .INP(n550), .ZN(n606) );
  XNOR3X1 U568 ( .IN1(keyinput96), .IN2(n542), .IN3(n607), .Q(N2768) );
  NAND2X0 U569 ( .IN1(keyinput105), .IN2(N46), .QN(n607) );
  AND3X1 U570 ( .IN1(n608), .IN2(n560), .IN3(n579), .Q(n542) );
  AND2X1 U571 ( .IN1(n524), .IN2(n521), .Q(n579) );
  XOR3X1 U572 ( .IN1(keyinput114), .IN2(n609), .IN3(n538), .Q(N2767) );
  NAND4X0 U573 ( .IN1(n523), .IN2(n608), .IN3(n590), .IN4(n591), .QN(n538) );
  NOR2X0 U574 ( .IN1(keyinput104), .IN2(n610), .QN(n609) );
  AO21X1 U575 ( .IN1(n611), .IN2(n612), .IN3(n613), .Q(N2762) );
  MUX21X1 U576 ( .IN1(n614), .IN2(n615), .S(keyinput109), .Q(n613) );
  NAND2X0 U577 ( .IN1(n616), .IN2(N28), .QN(n615) );
  XOR2X1 U578 ( .IN1(n547), .IN2(keyinput103), .Q(n616) );
  MUX21X1 U579 ( .IN1(n617), .IN2(n611), .S(keyinput103), .Q(n614) );
  NOR2X0 U580 ( .IN1(n611), .IN2(n612), .QN(n617) );
  INVX0 U581 ( .INP(n547), .ZN(n611) );
  NAND4X0 U582 ( .IN1(n521), .IN2(n608), .IN3(n525), .IN4(n560), .QN(n547) );
  NOR3X0 U583 ( .IN1(n514), .IN2(n584), .IN3(n510), .QN(n608) );
  INVX0 U584 ( .INP(n618), .ZN(n510) );
  AND2X1 U585 ( .IN1(n516), .IN2(n619), .Q(n584) );
  NAND3X0 U586 ( .IN1(n422), .IN2(n620), .IN3(N94), .QN(n619) );
  NOR2X0 U587 ( .IN1(n420), .IN2(N91), .QN(n422) );
  XOR3X1 U588 ( .IN1(keyinput110), .IN2(N10), .IN3(n532), .Q(N2756) );
  NAND4X0 U589 ( .IN1(n522), .IN2(n621), .IN3(n521), .IN4(n553), .QN(n532) );
  XOR2X1 U590 ( .IN1(n622), .IN2(n531), .Q(N2755) );
  NAND3X0 U591 ( .IN1(n525), .IN2(n621), .IN3(n554), .QN(n531) );
  XOR2X1 U592 ( .IN1(n623), .IN2(keyinput84), .Q(n525) );
  OR2X1 U593 ( .IN1(n590), .IN2(n624), .Q(n623) );
  XOR3X1 U594 ( .IN1(keyinput95), .IN2(N4), .IN3(n537), .Q(N2754) );
  NAND3X0 U595 ( .IN1(n621), .IN2(n524), .IN3(n554), .QN(n537) );
  NOR2X0 U596 ( .IN1(n560), .IN2(n521), .QN(n554) );
  INVX0 U597 ( .INP(n522), .ZN(n560) );
  AND2X1 U598 ( .IN1(n624), .IN2(n590), .Q(n524) );
  INVX0 U599 ( .INP(n591), .ZN(n624) );
  XOR2X1 U600 ( .IN1(n625), .IN2(n530), .Q(N2753) );
  NAND3X0 U601 ( .IN1(n523), .IN2(n553), .IN3(n621), .QN(n530) );
  AND2X1 U602 ( .IN1(n605), .IN2(n618), .Q(n621) );
  NOR2X0 U603 ( .IN1(n550), .IN2(n551), .QN(n618) );
  OA21X1 U604 ( .IN1(n566), .IN2(N76), .IN3(n626), .Q(n551) );
  XNOR2X1 U605 ( .IN1(n627), .IN2(keyinput87), .Q(n626) );
  NAND2X0 U606 ( .IN1(N76), .IN2(n566), .QN(n627) );
  AO21X1 U607 ( .IN1(n628), .IN2(n629), .IN3(N94), .Q(n566) );
  NAND2X0 U608 ( .IN1(n630), .IN2(n631), .QN(n629) );
  INVX0 U609 ( .INP(n632), .ZN(n630) );
  XOR2X1 U610 ( .IN1(n633), .IN2(keyinput80), .Q(n628) );
  NAND2X0 U611 ( .IN1(n634), .IN2(n632), .QN(n633) );
  NAND2X0 U612 ( .IN1(n635), .IN2(n636), .QN(n632) );
  XOR2X1 U613 ( .IN1(keyinput49), .IN2(n637), .Q(n636) );
  NOR2X0 U614 ( .IN1(n638), .IN2(n639), .QN(n637) );
  XOR2X1 U615 ( .IN1(keyinput27), .IN2(n481), .Q(n639) );
  XOR2X1 U616 ( .IN1(n640), .IN2(keyinput54), .Q(n635) );
  NAND2X0 U617 ( .IN1(n481), .IN2(n638), .QN(n640) );
  XNOR2X1 U618 ( .IN1(n641), .IN2(n482), .Q(n638) );
  NOR2X0 U619 ( .IN1(n642), .IN2(N40), .QN(n641) );
  INVX0 U620 ( .INP(keyinput14), .ZN(n642) );
  NOR2X0 U621 ( .IN1(n421), .IN2(N104), .QN(n481) );
  INVX0 U622 ( .INP(N66), .ZN(n421) );
  XOR2X1 U623 ( .IN1(keyinput78), .IN2(n631), .Q(n634) );
  MUX21X1 U624 ( .IN1(n480), .IN2(n643), .S(keyinput71), .Q(n631) );
  AOI21X1 U625 ( .IN1(n644), .IN2(n645), .IN3(n643), .QN(n480) );
  NOR2X0 U626 ( .IN1(n644), .IN2(n645), .QN(n643) );
  XNOR2X1 U627 ( .IN1(n646), .IN2(n436), .Q(n644) );
  XOR2X1 U628 ( .IN1(keyinput56), .IN2(n647), .Q(n436) );
  OA21X1 U629 ( .IN1(n648), .IN2(n612), .IN3(n649), .Q(n647) );
  XOR2X1 U630 ( .IN1(keyinput51), .IN2(n650), .Q(n649) );
  NOR2X0 U631 ( .IN1(N28), .IN2(n651), .QN(n650) );
  INVX0 U632 ( .INP(n651), .ZN(n648) );
  AO21X1 U633 ( .IN1(N43), .IN2(n652), .IN3(n653), .Q(n651) );
  XOR2X1 U634 ( .IN1(n654), .IN2(keyinput25), .Q(n653) );
  NAND2X0 U635 ( .IN1(n655), .IN2(n610), .QN(n654) );
  XOR2X1 U636 ( .IN1(n652), .IN2(keyinput13), .Q(n655) );
  AO21X1 U637 ( .IN1(n656), .IN2(n625), .IN3(n657), .Q(n646) );
  XOR2X1 U638 ( .IN1(keyinput44), .IN2(n658), .Q(n657) );
  NOR2X0 U639 ( .IN1(n659), .IN2(n660), .QN(n658) );
  XOR2X1 U640 ( .IN1(keyinput21), .IN2(N1), .Q(n660) );
  XOR2X1 U641 ( .IN1(keyinput45), .IN2(n659), .Q(n656) );
  XNOR2X1 U642 ( .IN1(n661), .IN2(keyinput38), .Q(n659) );
  OA21X1 U643 ( .IN1(n662), .IN2(N94), .IN3(N60), .Q(n550) );
  AOI21X1 U644 ( .IN1(n516), .IN2(n663), .IN3(n514), .QN(n605) );
  XNOR2X1 U645 ( .IN1(n664), .IN2(keyinput91), .Q(n514) );
  NAND2X0 U646 ( .IN1(n585), .IN2(n513), .QN(n664) );
  INVX0 U647 ( .INP(n575), .ZN(n513) );
  OA21X1 U648 ( .IN1(N72), .IN2(N94), .IN3(N53), .Q(n575) );
  XNOR2X1 U649 ( .IN1(keyinput88), .IN2(n665), .Q(n585) );
  OA21X1 U650 ( .IN1(n666), .IN2(n667), .IN3(n668), .Q(n665) );
  MUX21X1 U651 ( .IN1(n669), .IN2(n670), .S(n570), .Q(n668) );
  AND2X1 U652 ( .IN1(n671), .IN2(n489), .Q(n570) );
  XOR3X1 U653 ( .IN1(n672), .IN2(n496), .IN3(n487), .Q(n671) );
  XOR3X1 U654 ( .IN1(keyinput63), .IN2(n673), .IN3(n453), .Q(n487) );
  XOR3X1 U655 ( .IN1(keyinput30), .IN2(N22), .IN3(n482), .Q(n453) );
  OA21X1 U656 ( .IN1(n674), .IN2(n675), .IN3(n676), .Q(n673) );
  XOR2X1 U657 ( .IN1(keyinput62), .IN2(n677), .Q(n676) );
  NOR2X0 U658 ( .IN1(n457), .IN2(n455), .QN(n677) );
  INVX0 U659 ( .INP(n675), .ZN(n457) );
  AO21X1 U660 ( .IN1(n678), .IN2(n679), .IN3(n680), .Q(n675) );
  XOR2X1 U661 ( .IN1(keyinput46), .IN2(n681), .Q(n680) );
  NOR2X0 U662 ( .IN1(n679), .IN2(n678), .QN(n681) );
  INVX0 U663 ( .INP(n682), .ZN(n678) );
  MUX21X1 U664 ( .IN1(n683), .IN2(n684), .S(keyinput32), .Q(n682) );
  NAND2X0 U665 ( .IN1(N16), .IN2(n592), .QN(n683) );
  INVX0 U666 ( .INP(n455), .ZN(n674) );
  XOR3X1 U667 ( .IN1(keyinput39), .IN2(N1), .IN3(n661), .Q(n455) );
  XOR2X1 U668 ( .IN1(N4), .IN2(n622), .Q(n661) );
  XOR3X1 U669 ( .IN1(keyinput70), .IN2(N25), .IN3(n491), .Q(n672) );
  NOR2X0 U670 ( .IN1(n444), .IN2(N104), .QN(n491) );
  INVX0 U671 ( .INP(N63), .ZN(n444) );
  NAND2X0 U672 ( .IN1(n670), .IN2(n667), .QN(n669) );
  AND2X1 U673 ( .IN1(keyinput85), .IN2(n666), .Q(n670) );
  INVX0 U674 ( .INP(keyinput36), .ZN(n667) );
  INVX0 U675 ( .INP(n488), .ZN(n666) );
  OA21X1 U676 ( .IN1(N94), .IN2(N72), .IN3(N49), .Q(n488) );
  NAND4X0 U677 ( .IN1(N94), .IN2(N104), .IN3(n620), .IN4(n445), .QN(n663) );
  INVX0 U678 ( .INP(N88), .ZN(n445) );
  NAND3X0 U679 ( .IN1(n620), .IN2(n420), .IN3(N99), .QN(n516) );
  INVX0 U680 ( .INP(N104), .ZN(n420) );
  NAND2X0 U681 ( .IN1(N72), .IN2(N69), .QN(n620) );
  NOR2X0 U682 ( .IN1(n591), .IN2(n590), .QN(n553) );
  XOR2X1 U683 ( .IN1(keyinput79), .IN2(n685), .Q(n590) );
  AOI21X1 U684 ( .IN1(n577), .IN2(N82), .IN3(n574), .QN(n685) );
  NOR2X0 U685 ( .IN1(n577), .IN2(N82), .QN(n574) );
  NAND2X0 U686 ( .IN1(n469), .IN2(n489), .QN(n577) );
  XNOR3X1 U687 ( .IN1(n439), .IN2(n686), .IN3(n687), .Q(n469) );
  XNOR2X1 U688 ( .IN1(n688), .IN2(n689), .Q(n687) );
  OA21X1 U689 ( .IN1(n690), .IN2(n691), .IN3(keyinput61), .Q(n689) );
  XOR2X1 U690 ( .IN1(keyinput41), .IN2(n692), .Q(n691) );
  NOR2X0 U691 ( .IN1(N4), .IN2(n693), .QN(n692) );
  AND2X1 U692 ( .IN1(n693), .IN2(N4), .Q(n690) );
  AO21X1 U693 ( .IN1(N22), .IN2(n679), .IN3(n694), .Q(n693) );
  XOR2X1 U694 ( .IN1(n695), .IN2(keyinput19), .Q(n694) );
  OR2X1 U695 ( .IN1(n679), .IN2(N22), .Q(n695) );
  INVX0 U696 ( .INP(N13), .ZN(n679) );
  OA21X1 U697 ( .IN1(n696), .IN2(n697), .IN3(n698), .Q(n688) );
  MUX21X1 U698 ( .IN1(n699), .IN2(n700), .S(N46), .Q(n698) );
  NAND2X0 U699 ( .IN1(N43), .IN2(n696), .QN(n700) );
  XOR2X1 U700 ( .IN1(n610), .IN2(n696), .Q(n699) );
  NAND2X0 U701 ( .IN1(N53), .IN2(n701), .QN(n696) );
  XOR3X1 U702 ( .IN1(keyinput64), .IN2(N25), .IN3(n702), .Q(n686) );
  NOR2X0 U703 ( .IN1(N40), .IN2(keyinput16), .QN(n702) );
  AO21X1 U704 ( .IN1(n573), .IN2(n572), .IN3(n703), .Q(n591) );
  XOR2X1 U705 ( .IN1(n704), .IN2(keyinput74), .Q(n703) );
  OR2X1 U706 ( .IN1(n572), .IN2(n573), .Q(n704) );
  XOR2X1 U707 ( .IN1(N85), .IN2(keyinput4), .Q(n572) );
  NOR2X0 U708 ( .IN1(n464), .IN2(N94), .QN(n573) );
  XNOR2X1 U709 ( .IN1(n705), .IN2(n706), .Q(n464) );
  OA21X1 U710 ( .IN1(n707), .IN2(n708), .IN3(n709), .Q(n706) );
  XOR2X1 U711 ( .IN1(keyinput57), .IN2(n710), .Q(n709) );
  AND2X1 U712 ( .IN1(n708), .IN2(n707), .Q(n710) );
  AO21X1 U713 ( .IN1(n711), .IN2(n622), .IN3(n712), .Q(n708) );
  XOR2X1 U714 ( .IN1(keyinput40), .IN2(n713), .Q(n712) );
  NOR2X0 U715 ( .IN1(n622), .IN2(n711), .QN(n713) );
  INVX0 U716 ( .INP(N7), .ZN(n622) );
  XOR2X1 U717 ( .IN1(keyinput29), .IN2(n714), .Q(n711) );
  XOR2X1 U718 ( .IN1(N16), .IN2(n715), .Q(n714) );
  NOR2X0 U719 ( .IN1(N22), .IN2(keyinput17), .QN(n715) );
  INVX0 U720 ( .INP(n716), .ZN(n707) );
  MUX21X1 U721 ( .IN1(n717), .IN2(n718), .S(keyinput42), .Q(n716) );
  OA22X1 U722 ( .IN1(n437), .IN2(n719), .IN3(n720), .IN4(n721), .Q(n718) );
  XOR2X1 U723 ( .IN1(keyinput18), .IN2(N34), .Q(n721) );
  NAND2X0 U724 ( .IN1(n720), .IN2(n437), .QN(n717) );
  INVX0 U725 ( .INP(N34), .ZN(n437) );
  INVX0 U726 ( .INP(n719), .ZN(n720) );
  XNOR2X1 U727 ( .IN1(n612), .IN2(N43), .Q(n719) );
  NAND2X0 U728 ( .IN1(n722), .IN2(N56), .QN(n705) );
  XOR2X1 U729 ( .IN1(n723), .IN2(keyinput92), .Q(n523) );
  OR2X1 U730 ( .IN1(n521), .IN2(n522), .Q(n723) );
  XNOR2X1 U731 ( .IN1(N79), .IN2(n724), .Q(n522) );
  NOR2X0 U732 ( .IN1(N94), .IN2(n725), .QN(n724) );
  XOR2X1 U733 ( .IN1(keyinput81), .IN2(n726), .Q(n725) );
  OA21X1 U734 ( .IN1(n727), .IN2(n728), .IN3(n729), .Q(n726) );
  MUX21X1 U735 ( .IN1(n730), .IN2(n731), .S(n732), .Q(n729) );
  XOR2X1 U736 ( .IN1(keyinput43), .IN2(n733), .Q(n732) );
  OA21X1 U737 ( .IN1(n734), .IN2(n735), .IN3(n736), .Q(n733) );
  XOR2X1 U738 ( .IN1(keyinput31), .IN2(n737), .Q(n736) );
  NOR2X0 U739 ( .IN1(N1), .IN2(n406), .QN(n737) );
  INVX0 U740 ( .INP(n406), .ZN(n735) );
  XOR2X1 U741 ( .IN1(n738), .IN2(keyinput7), .Q(n406) );
  NAND2X0 U742 ( .IN1(N49), .IN2(n701), .QN(n738) );
  NOR2X0 U743 ( .IN1(N72), .IN2(N104), .QN(n701) );
  XOR2X1 U744 ( .IN1(n625), .IN2(keyinput8), .Q(n734) );
  NAND2X0 U745 ( .IN1(n730), .IN2(n728), .QN(n731) );
  AND2X1 U746 ( .IN1(keyinput53), .IN2(n727), .Q(n730) );
  INVX0 U747 ( .INP(keyinput77), .ZN(n728) );
  XOR3X1 U748 ( .IN1(keyinput75), .IN2(keyinput73), .IN3(n739), .Q(n727) );
  NAND2X0 U749 ( .IN1(n740), .IN2(n413), .QN(n739) );
  NAND2X0 U750 ( .IN1(n741), .IN2(n742), .QN(n413) );
  XNOR2X1 U751 ( .IN1(n411), .IN2(keyinput69), .Q(n740) );
  NOR2X0 U752 ( .IN1(n742), .IN2(n741), .QN(n411) );
  XNOR2X1 U753 ( .IN1(N13), .IN2(n684), .Q(n741) );
  XOR2X1 U754 ( .IN1(N16), .IN2(N19), .Q(n684) );
  XOR2X1 U755 ( .IN1(n645), .IN2(n496), .Q(n742) );
  XOR3X1 U756 ( .IN1(keyinput55), .IN2(N28), .IN3(n743), .Q(n496) );
  NAND2X0 U757 ( .IN1(n744), .IN2(n697), .QN(n743) );
  NAND2X0 U758 ( .IN1(N46), .IN2(n610), .QN(n697) );
  XOR2X1 U759 ( .IN1(n745), .IN2(keyinput33), .Q(n744) );
  NAND2X0 U760 ( .IN1(n746), .IN2(n652), .QN(n745) );
  XOR2X1 U761 ( .IN1(n610), .IN2(keyinput24), .Q(n746) );
  INVX0 U762 ( .INP(N43), .ZN(n610) );
  AO21X1 U763 ( .IN1(n439), .IN2(n747), .IN3(n748), .Q(n645) );
  XOR2X1 U764 ( .IN1(n749), .IN2(keyinput47), .Q(n748) );
  NAND2X0 U765 ( .IN1(n750), .IN2(n751), .QN(n749) );
  XNOR2X1 U766 ( .IN1(n439), .IN2(keyinput22), .Q(n750) );
  INVX0 U767 ( .INP(n751), .ZN(n747) );
  XOR2X1 U768 ( .IN1(n752), .IN2(N34), .Q(n751) );
  NAND2X0 U769 ( .IN1(keyinput26), .IN2(n438), .QN(n752) );
  XNOR2X1 U770 ( .IN1(n581), .IN2(keyinput1), .Q(n439) );
  INVX0 U771 ( .INP(N31), .ZN(n581) );
  XNOR2X1 U772 ( .IN1(n461), .IN2(n753), .Q(n521) );
  NOR2X0 U773 ( .IN1(n578), .IN2(keyinput37), .QN(n753) );
  AND2X1 U774 ( .IN1(n460), .IN2(n489), .Q(n578) );
  INVX0 U775 ( .INP(N94), .ZN(n489) );
  XNOR2X1 U776 ( .IN1(n754), .IN2(n755), .Q(n460) );
  XOR3X1 U777 ( .IN1(keyinput65), .IN2(keyinput34), .IN3(n756), .Q(n755) );
  OA21X1 U778 ( .IN1(n431), .IN2(n757), .IN3(n758), .Q(n756) );
  XOR2X1 U779 ( .IN1(n759), .IN2(keyinput52), .Q(n758) );
  NAND2X0 U780 ( .IN1(n431), .IN2(n652), .QN(n759) );
  INVX0 U781 ( .INP(N46), .ZN(n652) );
  XOR2X1 U782 ( .IN1(keyinput23), .IN2(N46), .Q(n757) );
  XOR2X1 U783 ( .IN1(n497), .IN2(N40), .Q(n431) );
  INVX0 U784 ( .INP(N25), .ZN(n497) );
  XOR3X1 U785 ( .IN1(n760), .IN2(n438), .IN3(n761), .Q(n754) );
  NAND2X0 U786 ( .IN1(n762), .IN2(keyinput58), .QN(n761) );
  XOR2X1 U787 ( .IN1(n482), .IN2(n763), .Q(n762) );
  OA21X1 U788 ( .IN1(N19), .IN2(n612), .IN3(n764), .Q(n763) );
  XOR2X1 U789 ( .IN1(keyinput20), .IN2(n765), .Q(n764) );
  NOR2X0 U790 ( .IN1(N28), .IN2(n592), .QN(n765) );
  INVX0 U791 ( .INP(N19), .ZN(n592) );
  INVX0 U792 ( .INP(N28), .ZN(n612) );
  XNOR2X1 U793 ( .IN1(N10), .IN2(keyinput0), .Q(n482) );
  XOR2X1 U794 ( .IN1(N37), .IN2(keyinput2), .Q(n438) );
  AND3X1 U795 ( .IN1(n722), .IN2(n766), .IN3(N60), .Q(n760) );
  INVX0 U796 ( .INP(keyinput9), .ZN(n766) );
  NOR2X0 U797 ( .IN1(n662), .IN2(N104), .QN(n722) );
  OA21X1 U798 ( .IN1(n662), .IN2(N94), .IN3(N56), .Q(n461) );
  INVX0 U799 ( .INP(N69), .ZN(n662) );
  INVX0 U800 ( .INP(N1), .ZN(n625) );
endmodule

