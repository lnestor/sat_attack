
module c6288 ( N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, 
        N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, 
        N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, N1901, 
        N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, 
        N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, 
        N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205,
         N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392,
         N409, N426, N443, N460, N477, N494, N511, N528, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241,
         N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180,
         N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280,
         N6287, N6288;
  wire   n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257;

  NAND2X0 U1675 ( .IN1(n1646), .IN2(n1647), .QN(N6288) );
  NAND3X0 U1676 ( .IN1(n1648), .IN2(n1649), .IN3(n1650), .QN(n1647) );
  AND2X1 U1677 ( .IN1(n1646), .IN2(n1651), .Q(N6287) );
  AO21X1 U1678 ( .IN1(n1648), .IN2(n1649), .IN3(n1650), .Q(n1646) );
  NAND2X0 U1679 ( .IN1(n1651), .IN2(n1652), .QN(n1650) );
  NAND4X0 U1680 ( .IN1(N528), .IN2(N256), .IN3(n1653), .IN4(n1654), .QN(n1652)
         );
  XOR2X1 U1681 ( .IN1(keyinput110), .IN2(n1655), .Q(n1651) );
  AOI22X1 U1682 ( .IN1(N256), .IN2(N528), .IN3(n1653), .IN4(n1656), .QN(n1655)
         );
  NAND2X0 U1683 ( .IN1(n1648), .IN2(n1657), .QN(N6280) );
  NAND3X0 U1684 ( .IN1(n1658), .IN2(n1659), .IN3(n1660), .QN(n1657) );
  AO21X1 U1685 ( .IN1(n1658), .IN2(n1659), .IN3(n1660), .Q(n1648) );
  NAND2X0 U1686 ( .IN1(n1649), .IN2(n1661), .QN(n1660) );
  NAND3X0 U1687 ( .IN1(n1662), .IN2(n1663), .IN3(n1664), .QN(n1661) );
  AO21X1 U1688 ( .IN1(n1664), .IN2(n1663), .IN3(n1662), .Q(n1649) );
  NAND2X0 U1689 ( .IN1(n1653), .IN2(n1665), .QN(n1662) );
  NAND3X0 U1690 ( .IN1(N239), .IN2(n1666), .IN3(N528), .QN(n1665) );
  AO21X1 U1691 ( .IN1(N528), .IN2(N239), .IN3(n1666), .Q(n1653) );
  NAND2X0 U1692 ( .IN1(n1667), .IN2(n1654), .QN(n1666) );
  OR2X1 U1693 ( .IN1(n1656), .IN2(N511), .Q(n1654) );
  MUX21X1 U1694 ( .IN1(n1656), .IN2(n1668), .S(N256), .Q(n1667) );
  NAND2X0 U1695 ( .IN1(N511), .IN2(n1656), .QN(n1668) );
  XOR2X1 U1696 ( .IN1(n1669), .IN2(keyinput104), .Q(n1656) );
  NAND2X0 U1697 ( .IN1(n1670), .IN2(n1671), .QN(n1669) );
  INVX0 U1698 ( .INP(n1672), .ZN(n1664) );
  NAND2X0 U1699 ( .IN1(n1658), .IN2(n1673), .QN(N6270) );
  NAND3X0 U1700 ( .IN1(n1674), .IN2(n1675), .IN3(n1676), .QN(n1673) );
  AO21X1 U1701 ( .IN1(n1674), .IN2(n1675), .IN3(n1676), .Q(n1658) );
  NAND2X0 U1702 ( .IN1(n1659), .IN2(n1677), .QN(n1676) );
  NAND3X0 U1703 ( .IN1(n1678), .IN2(n1679), .IN3(n1680), .QN(n1677) );
  AO21X1 U1704 ( .IN1(n1678), .IN2(n1679), .IN3(n1680), .Q(n1659) );
  AO21X1 U1705 ( .IN1(n1681), .IN2(n1682), .IN3(n1672), .Q(n1680) );
  XOR2X1 U1706 ( .IN1(n1683), .IN2(keyinput109), .Q(n1672) );
  OR2X1 U1707 ( .IN1(n1682), .IN2(n1681), .Q(n1683) );
  NAND2X0 U1708 ( .IN1(n1663), .IN2(n1684), .QN(n1682) );
  NAND3X0 U1709 ( .IN1(n1685), .IN2(n1686), .IN3(n1687), .QN(n1684) );
  AO21X1 U1710 ( .IN1(n1685), .IN2(n1686), .IN3(n1687), .Q(n1663) );
  AO21X1 U1711 ( .IN1(n1688), .IN2(n1689), .IN3(n1690), .Q(n1687) );
  INVX0 U1712 ( .INP(n1670), .ZN(n1690) );
  XOR2X1 U1713 ( .IN1(n1691), .IN2(keyinput102), .Q(n1670) );
  OR2X1 U1714 ( .IN1(n1689), .IN2(n1688), .Q(n1691) );
  NAND2X0 U1715 ( .IN1(n1671), .IN2(n1692), .QN(n1689) );
  NAND4X0 U1716 ( .IN1(N494), .IN2(N256), .IN3(n1693), .IN4(n1694), .QN(n1692)
         );
  AO22X1 U1717 ( .IN1(n1695), .IN2(n1693), .IN3(N494), .IN4(N256), .Q(n1671)
         );
  AND2X1 U1718 ( .IN1(N511), .IN2(N239), .Q(n1688) );
  AND2X1 U1719 ( .IN1(N222), .IN2(N528), .Q(n1681) );
  NAND2X0 U1720 ( .IN1(n1674), .IN2(n1696), .QN(N6260) );
  NAND3X0 U1721 ( .IN1(n1697), .IN2(n1698), .IN3(n1699), .QN(n1696) );
  AO21X1 U1722 ( .IN1(n1697), .IN2(n1698), .IN3(n1699), .Q(n1674) );
  NAND2X0 U1723 ( .IN1(n1675), .IN2(n1700), .QN(n1699) );
  NAND3X0 U1724 ( .IN1(n1701), .IN2(n1702), .IN3(n1703), .QN(n1700) );
  AO21X1 U1725 ( .IN1(n1701), .IN2(n1702), .IN3(n1703), .Q(n1675) );
  NAND2X0 U1726 ( .IN1(n1678), .IN2(n1704), .QN(n1703) );
  NAND3X0 U1727 ( .IN1(N528), .IN2(n1705), .IN3(N205), .QN(n1704) );
  AO21X1 U1728 ( .IN1(N205), .IN2(N528), .IN3(n1705), .Q(n1678) );
  NAND2X0 U1729 ( .IN1(n1679), .IN2(n1706), .QN(n1705) );
  NAND3X0 U1730 ( .IN1(n1707), .IN2(n1708), .IN3(n1709), .QN(n1706) );
  AO21X1 U1731 ( .IN1(n1707), .IN2(n1708), .IN3(n1709), .Q(n1679) );
  NAND2X0 U1732 ( .IN1(n1685), .IN2(n1710), .QN(n1709) );
  NAND3X0 U1733 ( .IN1(N511), .IN2(n1711), .IN3(N222), .QN(n1710) );
  AO21X1 U1734 ( .IN1(N222), .IN2(N511), .IN3(n1711), .Q(n1685) );
  NAND2X0 U1735 ( .IN1(n1686), .IN2(n1712), .QN(n1711) );
  NAND3X0 U1736 ( .IN1(n1713), .IN2(n1714), .IN3(n1715), .QN(n1712) );
  AO21X1 U1737 ( .IN1(n1713), .IN2(n1714), .IN3(n1715), .Q(n1686) );
  NAND2X0 U1738 ( .IN1(n1693), .IN2(n1716), .QN(n1715) );
  NAND3X0 U1739 ( .IN1(N494), .IN2(n1717), .IN3(N239), .QN(n1716) );
  AO21X1 U1740 ( .IN1(N239), .IN2(N494), .IN3(n1717), .Q(n1693) );
  NAND2X0 U1741 ( .IN1(n1718), .IN2(n1694), .QN(n1717) );
  OR2X1 U1742 ( .IN1(N477), .IN2(n1695), .Q(n1694) );
  MUX21X1 U1743 ( .IN1(n1695), .IN2(n1719), .S(N256), .Q(n1718) );
  NAND2X0 U1744 ( .IN1(n1695), .IN2(N477), .QN(n1719) );
  AOI21X1 U1745 ( .IN1(n1720), .IN2(n1721), .IN3(n1722), .QN(n1695) );
  INVX0 U1746 ( .INP(n1723), .ZN(n1722) );
  NAND2X0 U1747 ( .IN1(n1697), .IN2(n1724), .QN(N6250) );
  NAND3X0 U1748 ( .IN1(n1725), .IN2(n1726), .IN3(n1727), .QN(n1724) );
  AO21X1 U1749 ( .IN1(n1725), .IN2(n1726), .IN3(n1727), .Q(n1697) );
  NAND2X0 U1750 ( .IN1(n1698), .IN2(n1728), .QN(n1727) );
  NAND3X0 U1751 ( .IN1(n1729), .IN2(n1730), .IN3(n1731), .QN(n1728) );
  AO21X1 U1752 ( .IN1(n1729), .IN2(n1730), .IN3(n1731), .Q(n1698) );
  NAND2X0 U1753 ( .IN1(n1701), .IN2(n1732), .QN(n1731) );
  NAND3X0 U1754 ( .IN1(N528), .IN2(n1733), .IN3(N188), .QN(n1732) );
  AO21X1 U1755 ( .IN1(N188), .IN2(N528), .IN3(n1733), .Q(n1701) );
  NAND2X0 U1756 ( .IN1(n1702), .IN2(n1734), .QN(n1733) );
  NAND3X0 U1757 ( .IN1(n1735), .IN2(n1736), .IN3(n1737), .QN(n1734) );
  AO21X1 U1758 ( .IN1(n1735), .IN2(n1736), .IN3(n1737), .Q(n1702) );
  NAND2X0 U1759 ( .IN1(n1707), .IN2(n1738), .QN(n1737) );
  NAND3X0 U1760 ( .IN1(N511), .IN2(n1739), .IN3(N205), .QN(n1738) );
  AO21X1 U1761 ( .IN1(N205), .IN2(N511), .IN3(n1739), .Q(n1707) );
  NAND2X0 U1762 ( .IN1(n1708), .IN2(n1740), .QN(n1739) );
  NAND3X0 U1763 ( .IN1(n1741), .IN2(n1742), .IN3(n1743), .QN(n1740) );
  AO21X1 U1764 ( .IN1(n1741), .IN2(n1742), .IN3(n1743), .Q(n1708) );
  NAND2X0 U1765 ( .IN1(n1713), .IN2(n1744), .QN(n1743) );
  NAND3X0 U1766 ( .IN1(N494), .IN2(n1745), .IN3(N222), .QN(n1744) );
  AO21X1 U1767 ( .IN1(N222), .IN2(N494), .IN3(n1745), .Q(n1713) );
  NAND2X0 U1768 ( .IN1(n1714), .IN2(n1746), .QN(n1745) );
  NAND3X0 U1769 ( .IN1(n1747), .IN2(n1748), .IN3(n1749), .QN(n1746) );
  AO21X1 U1770 ( .IN1(n1747), .IN2(n1748), .IN3(n1749), .Q(n1714) );
  NAND2X0 U1771 ( .IN1(n1723), .IN2(n1750), .QN(n1749) );
  NAND3X0 U1772 ( .IN1(N477), .IN2(N239), .IN3(n1751), .QN(n1750) );
  AO21X1 U1773 ( .IN1(N477), .IN2(N239), .IN3(n1751), .Q(n1723) );
  XNOR2X1 U1774 ( .IN1(n1721), .IN2(n1720), .Q(n1751) );
  NAND2X0 U1775 ( .IN1(N460), .IN2(N256), .QN(n1720) );
  AO21X1 U1776 ( .IN1(n1752), .IN2(n1753), .IN3(n1754), .Q(n1721) );
  INVX0 U1777 ( .INP(n1755), .ZN(n1754) );
  NAND2X0 U1778 ( .IN1(n1725), .IN2(n1756), .QN(N6240) );
  NAND3X0 U1779 ( .IN1(n1757), .IN2(n1758), .IN3(n1759), .QN(n1756) );
  AO21X1 U1780 ( .IN1(n1757), .IN2(n1758), .IN3(n1759), .Q(n1725) );
  NAND2X0 U1781 ( .IN1(n1726), .IN2(n1760), .QN(n1759) );
  NAND3X0 U1782 ( .IN1(n1761), .IN2(n1762), .IN3(n1763), .QN(n1760) );
  AO21X1 U1783 ( .IN1(n1761), .IN2(n1762), .IN3(n1763), .Q(n1726) );
  NAND2X0 U1784 ( .IN1(n1729), .IN2(n1764), .QN(n1763) );
  NAND3X0 U1785 ( .IN1(N528), .IN2(n1765), .IN3(N171), .QN(n1764) );
  AO21X1 U1786 ( .IN1(N171), .IN2(N528), .IN3(n1765), .Q(n1729) );
  NAND2X0 U1787 ( .IN1(n1730), .IN2(n1766), .QN(n1765) );
  NAND3X0 U1788 ( .IN1(n1767), .IN2(n1768), .IN3(n1769), .QN(n1766) );
  AO21X1 U1789 ( .IN1(n1767), .IN2(n1768), .IN3(n1769), .Q(n1730) );
  NAND2X0 U1790 ( .IN1(n1735), .IN2(n1770), .QN(n1769) );
  NAND3X0 U1791 ( .IN1(N511), .IN2(n1771), .IN3(N188), .QN(n1770) );
  AO21X1 U1792 ( .IN1(N188), .IN2(N511), .IN3(n1771), .Q(n1735) );
  NAND2X0 U1793 ( .IN1(n1736), .IN2(n1772), .QN(n1771) );
  NAND3X0 U1794 ( .IN1(n1773), .IN2(n1774), .IN3(n1775), .QN(n1772) );
  AO21X1 U1795 ( .IN1(n1773), .IN2(n1774), .IN3(n1775), .Q(n1736) );
  XOR2X1 U1796 ( .IN1(n1776), .IN2(keyinput100), .Q(n1775) );
  NAND2X0 U1797 ( .IN1(n1741), .IN2(n1777), .QN(n1776) );
  NAND3X0 U1798 ( .IN1(N494), .IN2(n1778), .IN3(N205), .QN(n1777) );
  AO21X1 U1799 ( .IN1(N205), .IN2(N494), .IN3(n1778), .Q(n1741) );
  NAND2X0 U1800 ( .IN1(n1742), .IN2(n1779), .QN(n1778) );
  NAND3X0 U1801 ( .IN1(n1780), .IN2(n1781), .IN3(n1782), .QN(n1779) );
  AO21X1 U1802 ( .IN1(n1780), .IN2(n1781), .IN3(n1782), .Q(n1742) );
  NAND2X0 U1803 ( .IN1(n1747), .IN2(n1783), .QN(n1782) );
  NAND3X0 U1804 ( .IN1(N477), .IN2(n1784), .IN3(N222), .QN(n1783) );
  AO21X1 U1805 ( .IN1(N222), .IN2(N477), .IN3(n1784), .Q(n1747) );
  NAND2X0 U1806 ( .IN1(n1748), .IN2(n1785), .QN(n1784) );
  NAND3X0 U1807 ( .IN1(n1786), .IN2(n1787), .IN3(n1788), .QN(n1785) );
  AO21X1 U1808 ( .IN1(n1786), .IN2(n1787), .IN3(n1788), .Q(n1748) );
  NAND2X0 U1809 ( .IN1(n1755), .IN2(n1789), .QN(n1788) );
  NAND3X0 U1810 ( .IN1(N460), .IN2(N239), .IN3(n1790), .QN(n1789) );
  AO21X1 U1811 ( .IN1(N460), .IN2(N239), .IN3(n1790), .Q(n1755) );
  XNOR2X1 U1812 ( .IN1(n1753), .IN2(n1752), .Q(n1790) );
  XNOR2X1 U1813 ( .IN1(keyinput82), .IN2(n1791), .Q(n1752) );
  OA21X1 U1814 ( .IN1(n1792), .IN2(n1793), .IN3(n1794), .Q(n1791) );
  NAND2X0 U1815 ( .IN1(N443), .IN2(N256), .QN(n1753) );
  INVX0 U1816 ( .INP(n1795), .ZN(n1781) );
  NAND2X0 U1817 ( .IN1(n1757), .IN2(n1796), .QN(N6230) );
  NAND3X0 U1818 ( .IN1(n1797), .IN2(n1798), .IN3(n1799), .QN(n1796) );
  AO21X1 U1819 ( .IN1(n1797), .IN2(n1798), .IN3(n1799), .Q(n1757) );
  NAND2X0 U1820 ( .IN1(n1758), .IN2(n1800), .QN(n1799) );
  NAND3X0 U1821 ( .IN1(n1801), .IN2(n1802), .IN3(n1803), .QN(n1800) );
  AO21X1 U1822 ( .IN1(n1803), .IN2(n1802), .IN3(n1801), .Q(n1758) );
  NAND2X0 U1823 ( .IN1(n1761), .IN2(n1804), .QN(n1801) );
  NAND3X0 U1824 ( .IN1(N154), .IN2(N528), .IN3(n1805), .QN(n1804) );
  AO21X1 U1825 ( .IN1(N154), .IN2(N528), .IN3(n1805), .Q(n1761) );
  XOR2X1 U1826 ( .IN1(n1806), .IN2(keyinput115), .Q(n1805) );
  NAND2X0 U1827 ( .IN1(n1762), .IN2(n1807), .QN(n1806) );
  NAND3X0 U1828 ( .IN1(n1808), .IN2(n1809), .IN3(n1810), .QN(n1807) );
  AO21X1 U1829 ( .IN1(n1810), .IN2(n1809), .IN3(n1808), .Q(n1762) );
  NAND2X0 U1830 ( .IN1(n1767), .IN2(n1811), .QN(n1808) );
  NAND3X0 U1831 ( .IN1(N511), .IN2(n1812), .IN3(N171), .QN(n1811) );
  AO21X1 U1832 ( .IN1(N171), .IN2(N511), .IN3(n1812), .Q(n1767) );
  NAND2X0 U1833 ( .IN1(n1768), .IN2(n1813), .QN(n1812) );
  NAND3X0 U1834 ( .IN1(n1814), .IN2(n1815), .IN3(n1816), .QN(n1813) );
  AO21X1 U1835 ( .IN1(n1814), .IN2(n1815), .IN3(n1816), .Q(n1768) );
  NAND2X0 U1836 ( .IN1(n1773), .IN2(n1817), .QN(n1816) );
  NAND3X0 U1837 ( .IN1(N494), .IN2(n1818), .IN3(N188), .QN(n1817) );
  AO21X1 U1838 ( .IN1(N188), .IN2(N494), .IN3(n1818), .Q(n1773) );
  NAND2X0 U1839 ( .IN1(n1774), .IN2(n1819), .QN(n1818) );
  NAND3X0 U1840 ( .IN1(n1820), .IN2(n1821), .IN3(n1822), .QN(n1819) );
  AO21X1 U1841 ( .IN1(n1822), .IN2(n1821), .IN3(n1820), .Q(n1774) );
  AO21X1 U1842 ( .IN1(n1823), .IN2(n1824), .IN3(n1795), .Q(n1820) );
  NOR2X0 U1843 ( .IN1(n1824), .IN2(n1823), .QN(n1795) );
  XOR2X1 U1844 ( .IN1(n1825), .IN2(keyinput20), .Q(n1824) );
  NAND2X0 U1845 ( .IN1(N205), .IN2(N477), .QN(n1825) );
  AOI21X1 U1846 ( .IN1(n1826), .IN2(n1780), .IN3(n1827), .QN(n1823) );
  XOR2X1 U1847 ( .IN1(keyinput94), .IN2(n1828), .Q(n1827) );
  AOI21X1 U1848 ( .IN1(n1829), .IN2(n1830), .IN3(n1831), .QN(n1828) );
  INVX0 U1849 ( .INP(n1780), .ZN(n1831) );
  AO21X1 U1850 ( .IN1(n1830), .IN2(n1829), .IN3(n1832), .Q(n1780) );
  XNOR2X1 U1851 ( .IN1(keyinput91), .IN2(n1833), .Q(n1832) );
  XOR2X1 U1852 ( .IN1(n1833), .IN2(keyinput91), .Q(n1826) );
  NAND2X0 U1853 ( .IN1(n1786), .IN2(n1834), .QN(n1833) );
  NAND3X0 U1854 ( .IN1(N460), .IN2(n1835), .IN3(N222), .QN(n1834) );
  AO21X1 U1855 ( .IN1(N222), .IN2(N460), .IN3(n1835), .Q(n1786) );
  NAND2X0 U1856 ( .IN1(n1787), .IN2(n1836), .QN(n1835) );
  NAND3X0 U1857 ( .IN1(n1837), .IN2(n1838), .IN3(n1839), .QN(n1836) );
  AO21X1 U1858 ( .IN1(n1837), .IN2(n1838), .IN3(n1839), .Q(n1787) );
  XNOR2X1 U1859 ( .IN1(n1792), .IN2(n1793), .Q(n1839) );
  NAND2X0 U1860 ( .IN1(n1794), .IN2(n1840), .QN(n1793) );
  NAND4X0 U1861 ( .IN1(N426), .IN2(N256), .IN3(n1841), .IN4(n1842), .QN(n1840)
         );
  AO22X1 U1862 ( .IN1(n1843), .IN2(n1841), .IN3(N426), .IN4(N256), .Q(n1794)
         );
  AND2X1 U1863 ( .IN1(N239), .IN2(N443), .Q(n1792) );
  INVX0 U1864 ( .INP(n1844), .ZN(n1838) );
  INVX0 U1865 ( .INP(n1845), .ZN(n1822) );
  INVX0 U1866 ( .INP(n1846), .ZN(n1803) );
  NAND2X0 U1867 ( .IN1(n1797), .IN2(n1847), .QN(N6220) );
  NAND3X0 U1868 ( .IN1(n1848), .IN2(n1849), .IN3(n1850), .QN(n1847) );
  AO21X1 U1869 ( .IN1(n1848), .IN2(n1849), .IN3(n1850), .Q(n1797) );
  OAI21X1 U1870 ( .IN1(n1851), .IN2(n1852), .IN3(n1798), .QN(n1850) );
  NAND2X0 U1871 ( .IN1(n1853), .IN2(n1851), .QN(n1798) );
  XOR2X1 U1872 ( .IN1(n1854), .IN2(n1855), .Q(n1853) );
  AOI21X1 U1873 ( .IN1(n1855), .IN2(n1854), .IN3(n1846), .QN(n1852) );
  NOR2X0 U1874 ( .IN1(n1854), .IN2(n1855), .QN(n1846) );
  NAND2X0 U1875 ( .IN1(n1802), .IN2(n1856), .QN(n1854) );
  NAND3X0 U1876 ( .IN1(n1857), .IN2(n1858), .IN3(n1859), .QN(n1856) );
  AO21X1 U1877 ( .IN1(n1857), .IN2(n1858), .IN3(n1859), .Q(n1802) );
  AO21X1 U1878 ( .IN1(n1860), .IN2(n1861), .IN3(n1862), .Q(n1859) );
  INVX0 U1879 ( .INP(n1810), .ZN(n1862) );
  XOR2X1 U1880 ( .IN1(n1863), .IN2(keyinput108), .Q(n1810) );
  OR2X1 U1881 ( .IN1(n1861), .IN2(n1860), .Q(n1863) );
  AND2X1 U1882 ( .IN1(n1864), .IN2(n1865), .Q(n1861) );
  NAND3X0 U1883 ( .IN1(n1866), .IN2(n1814), .IN3(n1809), .QN(n1865) );
  XNOR2X1 U1884 ( .IN1(keyinput107), .IN2(n1867), .Q(n1864) );
  OA21X1 U1885 ( .IN1(n1868), .IN2(n1869), .IN3(n1809), .Q(n1867) );
  NAND3X0 U1886 ( .IN1(n1866), .IN2(n1814), .IN3(n1870), .QN(n1809) );
  OR2X1 U1887 ( .IN1(n1869), .IN2(n1868), .Q(n1870) );
  AO21X1 U1888 ( .IN1(N171), .IN2(N494), .IN3(n1871), .Q(n1814) );
  NAND3X0 U1889 ( .IN1(N494), .IN2(n1871), .IN3(N171), .QN(n1866) );
  NAND2X0 U1890 ( .IN1(n1815), .IN2(n1872), .QN(n1871) );
  NAND3X0 U1891 ( .IN1(n1873), .IN2(n1874), .IN3(n1875), .QN(n1872) );
  AO21X1 U1892 ( .IN1(n1873), .IN2(n1874), .IN3(n1875), .Q(n1815) );
  AO21X1 U1893 ( .IN1(n1876), .IN2(n1877), .IN3(n1845), .Q(n1875) );
  NOR2X0 U1894 ( .IN1(n1877), .IN2(n1876), .QN(n1845) );
  NAND2X0 U1895 ( .IN1(n1821), .IN2(n1878), .QN(n1877) );
  NAND3X0 U1896 ( .IN1(n1879), .IN2(n1880), .IN3(n1881), .QN(n1878) );
  AO21X1 U1897 ( .IN1(n1879), .IN2(n1880), .IN3(n1881), .Q(n1821) );
  XNOR2X1 U1898 ( .IN1(n1882), .IN2(keyinput93), .Q(n1881) );
  NAND2X0 U1899 ( .IN1(n1830), .IN2(n1883), .QN(n1882) );
  NAND3X0 U1900 ( .IN1(N460), .IN2(n1884), .IN3(N205), .QN(n1883) );
  AO21X1 U1901 ( .IN1(N205), .IN2(N460), .IN3(n1884), .Q(n1830) );
  NAND2X0 U1902 ( .IN1(n1829), .IN2(n1885), .QN(n1884) );
  NAND3X0 U1903 ( .IN1(n1886), .IN2(n1887), .IN3(n1888), .QN(n1885) );
  AO21X1 U1904 ( .IN1(n1886), .IN2(n1887), .IN3(n1888), .Q(n1829) );
  NAND2X0 U1905 ( .IN1(n1837), .IN2(n1889), .QN(n1888) );
  NAND3X0 U1906 ( .IN1(N443), .IN2(n1890), .IN3(N222), .QN(n1889) );
  AO21X1 U1907 ( .IN1(N222), .IN2(N443), .IN3(n1890), .Q(n1837) );
  AO21X1 U1908 ( .IN1(n1891), .IN2(n1892), .IN3(n1844), .Q(n1890) );
  NOR2X0 U1909 ( .IN1(n1892), .IN2(n1891), .QN(n1844) );
  NAND2X0 U1910 ( .IN1(n1841), .IN2(n1893), .QN(n1892) );
  NAND3X0 U1911 ( .IN1(N239), .IN2(n1894), .IN3(N426), .QN(n1893) );
  AO21X1 U1912 ( .IN1(N426), .IN2(N239), .IN3(n1894), .Q(n1841) );
  NAND2X0 U1913 ( .IN1(n1895), .IN2(n1842), .QN(n1894) );
  OR2X1 U1914 ( .IN1(N409), .IN2(n1843), .Q(n1842) );
  MUX21X1 U1915 ( .IN1(n1843), .IN2(n1896), .S(N256), .Q(n1895) );
  NAND2X0 U1916 ( .IN1(n1843), .IN2(N409), .QN(n1896) );
  OA21X1 U1917 ( .IN1(n1897), .IN2(n1898), .IN3(n1899), .Q(n1843) );
  XNOR2X1 U1918 ( .IN1(keyinput74), .IN2(n1900), .Q(n1891) );
  OA21X1 U1919 ( .IN1(n1901), .IN2(n1902), .IN3(n1903), .Q(n1900) );
  INVX0 U1920 ( .INP(n1904), .ZN(n1880) );
  XNOR2X1 U1921 ( .IN1(n1905), .IN2(keyinput18), .Q(n1876) );
  NAND2X0 U1922 ( .IN1(N188), .IN2(N477), .QN(n1905) );
  INVX0 U1923 ( .INP(n1906), .ZN(n1868) );
  NOR2X0 U1924 ( .IN1(n1907), .IN2(n1908), .QN(n1860) );
  XOR2X1 U1925 ( .IN1(n1909), .IN2(keyinput14), .Q(n1855) );
  NAND2X0 U1926 ( .IN1(N137), .IN2(N528), .QN(n1909) );
  XNOR2X1 U1927 ( .IN1(n1910), .IN2(keyinput121), .Q(n1851) );
  NAND2X0 U1928 ( .IN1(n1911), .IN2(n1912), .QN(n1910) );
  INVX0 U1929 ( .INP(n1913), .ZN(n1912) );
  NOR2X0 U1930 ( .IN1(n1914), .IN2(n1915), .QN(N6210) );
  XOR2X1 U1931 ( .IN1(keyinput127), .IN2(n1916), .Q(n1915) );
  NOR2X0 U1932 ( .IN1(n1917), .IN2(n1918), .QN(n1916) );
  AOI21X1 U1933 ( .IN1(n1919), .IN2(n1920), .IN3(n1917), .QN(n1914) );
  INVX0 U1934 ( .INP(n1848), .ZN(n1917) );
  AO21X1 U1935 ( .IN1(n1920), .IN2(n1919), .IN3(n1918), .Q(n1848) );
  XOR2X1 U1936 ( .IN1(n1921), .IN2(keyinput123), .Q(n1918) );
  NAND2X0 U1937 ( .IN1(n1849), .IN2(n1922), .QN(n1921) );
  NAND3X0 U1938 ( .IN1(n1923), .IN2(n1924), .IN3(n1925), .QN(n1922) );
  AO21X1 U1939 ( .IN1(n1923), .IN2(n1924), .IN3(n1925), .Q(n1849) );
  AO21X1 U1940 ( .IN1(n1926), .IN2(n1927), .IN3(n1913), .Q(n1925) );
  NOR2X0 U1941 ( .IN1(n1927), .IN2(n1926), .QN(n1913) );
  NAND2X0 U1942 ( .IN1(n1911), .IN2(n1928), .QN(n1927) );
  NAND3X0 U1943 ( .IN1(n1929), .IN2(n1930), .IN3(n1931), .QN(n1928) );
  AO21X1 U1944 ( .IN1(n1929), .IN2(n1930), .IN3(n1931), .Q(n1911) );
  XNOR2X1 U1945 ( .IN1(n1932), .IN2(keyinput114), .Q(n1931) );
  NAND2X0 U1946 ( .IN1(n1857), .IN2(n1933), .QN(n1932) );
  NAND3X0 U1947 ( .IN1(N511), .IN2(n1934), .IN3(N137), .QN(n1933) );
  AO21X1 U1948 ( .IN1(N137), .IN2(N511), .IN3(n1934), .Q(n1857) );
  NAND2X0 U1949 ( .IN1(n1858), .IN2(n1935), .QN(n1934) );
  NAND3X0 U1950 ( .IN1(n1936), .IN2(n1937), .IN3(n1938), .QN(n1935) );
  AO21X1 U1951 ( .IN1(n1938), .IN2(n1937), .IN3(n1936), .Q(n1858) );
  AO21X1 U1952 ( .IN1(n1939), .IN2(n1940), .IN3(n1869), .Q(n1936) );
  XOR2X1 U1953 ( .IN1(n1941), .IN2(keyinput101), .Q(n1869) );
  OR2X1 U1954 ( .IN1(n1940), .IN2(n1939), .Q(n1941) );
  NAND2X0 U1955 ( .IN1(n1906), .IN2(n1942), .QN(n1940) );
  NAND3X0 U1956 ( .IN1(n1943), .IN2(n1944), .IN3(n1945), .QN(n1942) );
  AO21X1 U1957 ( .IN1(n1943), .IN2(n1944), .IN3(n1945), .Q(n1906) );
  NAND2X0 U1958 ( .IN1(n1873), .IN2(n1946), .QN(n1945) );
  NAND4X0 U1959 ( .IN1(N171), .IN2(N477), .IN3(n1947), .IN4(n1948), .QN(n1946)
         );
  AO22X1 U1960 ( .IN1(N171), .IN2(N477), .IN3(n1947), .IN4(n1948), .Q(n1873)
         );
  NAND2X0 U1961 ( .IN1(n1949), .IN2(n1874), .QN(n1948) );
  XOR2X1 U1962 ( .IN1(keyinput96), .IN2(n1950), .Q(n1947) );
  OA21X1 U1963 ( .IN1(n1951), .IN2(n1952), .IN3(n1874), .Q(n1950) );
  OAI21X1 U1964 ( .IN1(n1952), .IN2(n1951), .IN3(n1949), .QN(n1874) );
  AOI21X1 U1965 ( .IN1(n1953), .IN2(n1954), .IN3(n1904), .QN(n1949) );
  NOR2X0 U1966 ( .IN1(n1954), .IN2(n1953), .QN(n1904) );
  NAND2X0 U1967 ( .IN1(n1879), .IN2(n1955), .QN(n1954) );
  NAND3X0 U1968 ( .IN1(n1956), .IN2(n1957), .IN3(n1958), .QN(n1955) );
  AO21X1 U1969 ( .IN1(n1956), .IN2(n1957), .IN3(n1958), .Q(n1879) );
  NAND2X0 U1970 ( .IN1(n1886), .IN2(n1959), .QN(n1958) );
  NAND3X0 U1971 ( .IN1(N443), .IN2(n1960), .IN3(N205), .QN(n1959) );
  AO21X1 U1972 ( .IN1(N205), .IN2(N443), .IN3(n1960), .Q(n1886) );
  NAND2X0 U1973 ( .IN1(n1887), .IN2(n1961), .QN(n1960) );
  NAND3X0 U1974 ( .IN1(n1962), .IN2(n1963), .IN3(n1964), .QN(n1961) );
  AO21X1 U1975 ( .IN1(n1964), .IN2(n1962), .IN3(n1963), .Q(n1887) );
  XNOR2X1 U1976 ( .IN1(n1901), .IN2(n1902), .Q(n1963) );
  AND2X1 U1977 ( .IN1(N222), .IN2(N426), .Q(n1902) );
  NAND2X0 U1978 ( .IN1(n1903), .IN2(n1965), .QN(n1901) );
  NAND3X0 U1979 ( .IN1(n1966), .IN2(n1967), .IN3(n1968), .QN(n1965) );
  AO21X1 U1980 ( .IN1(n1966), .IN2(n1967), .IN3(n1968), .Q(n1903) );
  NAND2X0 U1981 ( .IN1(n1899), .IN2(n1969), .QN(n1968) );
  NAND3X0 U1982 ( .IN1(N239), .IN2(n1970), .IN3(N409), .QN(n1969) );
  AO21X1 U1983 ( .IN1(N409), .IN2(N239), .IN3(n1970), .Q(n1899) );
  XOR3X1 U1984 ( .IN1(keyinput60), .IN2(n1897), .IN3(n1898), .Q(n1970) );
  AOI22X1 U1985 ( .IN1(n1971), .IN2(n1972), .IN3(n1973), .IN4(n1974), .QN(
        n1898) );
  NOR2X0 U1986 ( .IN1(n1975), .IN2(n1976), .QN(n1897) );
  XOR2X1 U1987 ( .IN1(n1977), .IN2(keyinput17), .Q(n1953) );
  NAND2X0 U1988 ( .IN1(N188), .IN2(N460), .QN(n1977) );
  INVX0 U1989 ( .INP(n1978), .ZN(n1951) );
  AND2X1 U1990 ( .IN1(N154), .IN2(N494), .Q(n1939) );
  INVX0 U1991 ( .INP(n1979), .ZN(n1938) );
  XOR2X1 U1992 ( .IN1(n1980), .IN2(keyinput12), .Q(n1926) );
  NAND2X0 U1993 ( .IN1(N120), .IN2(N528), .QN(n1980) );
  NAND2X0 U1994 ( .IN1(n1920), .IN2(n1981), .QN(N6200) );
  NAND3X0 U1995 ( .IN1(n1982), .IN2(n1983), .IN3(n1984), .QN(n1981) );
  AO21X1 U1996 ( .IN1(n1982), .IN2(n1983), .IN3(n1984), .Q(n1920) );
  NAND2X0 U1997 ( .IN1(n1919), .IN2(n1985), .QN(n1984) );
  AO221X1 U1998 ( .IN1(n1986), .IN2(n1923), .IN3(n1987), .IN4(n1988), .IN5(
        n1989), .Q(n1985) );
  NAND3X0 U1999 ( .IN1(n1986), .IN2(n1923), .IN3(n1990), .QN(n1919) );
  AO21X1 U2000 ( .IN1(n1987), .IN2(n1988), .IN3(n1989), .Q(n1990) );
  AO21X1 U2001 ( .IN1(N103), .IN2(N528), .IN3(n1991), .Q(n1923) );
  NAND3X0 U2002 ( .IN1(N528), .IN2(n1991), .IN3(N103), .QN(n1986) );
  NAND2X0 U2003 ( .IN1(n1924), .IN2(n1992), .QN(n1991) );
  NAND4X0 U2004 ( .IN1(n1993), .IN2(n1994), .IN3(n1995), .IN4(n1996), .QN(
        n1992) );
  AO22X1 U2005 ( .IN1(n1995), .IN2(n1996), .IN3(n1993), .IN4(n1994), .Q(n1924)
         );
  AO21X1 U2006 ( .IN1(N120), .IN2(N511), .IN3(n1997), .Q(n1994) );
  XNOR2X1 U2007 ( .IN1(n1998), .IN2(keyinput113), .Q(n1993) );
  NAND2X0 U2008 ( .IN1(n1999), .IN2(n1929), .QN(n1998) );
  INVX0 U2009 ( .INP(n1997), .ZN(n1929) );
  OA21X1 U2010 ( .IN1(n2000), .IN2(n1908), .IN3(n1999), .Q(n1997) );
  AND2X1 U2011 ( .IN1(n1930), .IN2(n2001), .Q(n1999) );
  NAND3X0 U2012 ( .IN1(n2002), .IN2(n2003), .IN3(n2004), .QN(n2001) );
  AO21X1 U2013 ( .IN1(n2002), .IN2(n2003), .IN3(n2004), .Q(n1930) );
  AO21X1 U2014 ( .IN1(n2005), .IN2(n2006), .IN3(n1979), .Q(n2004) );
  XOR2X1 U2015 ( .IN1(n2007), .IN2(keyinput103), .Q(n1979) );
  OR2X1 U2016 ( .IN1(n2006), .IN2(n2005), .Q(n2007) );
  NAND2X0 U2017 ( .IN1(n1937), .IN2(n2008), .QN(n2006) );
  NAND3X0 U2018 ( .IN1(n2009), .IN2(n2010), .IN3(n2011), .QN(n2008) );
  AO21X1 U2019 ( .IN1(n2009), .IN2(n2010), .IN3(n2011), .Q(n1937) );
  NAND2X0 U2020 ( .IN1(n1943), .IN2(n2012), .QN(n2011) );
  NAND3X0 U2021 ( .IN1(N477), .IN2(n2013), .IN3(N154), .QN(n2012) );
  AO21X1 U2022 ( .IN1(N154), .IN2(N477), .IN3(n2013), .Q(n1943) );
  NAND2X0 U2023 ( .IN1(n1944), .IN2(n2014), .QN(n2013) );
  NAND3X0 U2024 ( .IN1(n2015), .IN2(n2016), .IN3(n2017), .QN(n2014) );
  AO21X1 U2025 ( .IN1(n2015), .IN2(n2016), .IN3(n2017), .Q(n1944) );
  AO21X1 U2026 ( .IN1(n2018), .IN2(n2019), .IN3(n1952), .Q(n2017) );
  XNOR2X1 U2027 ( .IN1(n2020), .IN2(keyinput92), .Q(n1952) );
  OR2X1 U2028 ( .IN1(n2019), .IN2(n2018), .Q(n2020) );
  NAND2X0 U2029 ( .IN1(n1978), .IN2(n2021), .QN(n2019) );
  NAND3X0 U2030 ( .IN1(n2022), .IN2(n2023), .IN3(n2024), .QN(n2021) );
  AO21X1 U2031 ( .IN1(n2022), .IN2(n2023), .IN3(n2024), .Q(n1978) );
  NAND2X0 U2032 ( .IN1(n1956), .IN2(n2025), .QN(n2024) );
  NAND3X0 U2033 ( .IN1(N443), .IN2(n2026), .IN3(N188), .QN(n2025) );
  AO21X1 U2034 ( .IN1(N188), .IN2(N443), .IN3(n2026), .Q(n1956) );
  XOR2X1 U2035 ( .IN1(keyinput84), .IN2(n2027), .Q(n2026) );
  NOR2X0 U2036 ( .IN1(n2028), .IN2(n2029), .QN(n2027) );
  XOR2X1 U2037 ( .IN1(n2030), .IN2(keyinput81), .Q(n2029) );
  NAND2X0 U2038 ( .IN1(n2031), .IN2(n1957), .QN(n2030) );
  OA21X1 U2039 ( .IN1(n2032), .IN2(n2033), .IN3(n1957), .Q(n2028) );
  OAI21X1 U2040 ( .IN1(n2032), .IN2(n2033), .IN3(n2031), .QN(n1957) );
  AOI21X1 U2041 ( .IN1(n2034), .IN2(n2035), .IN3(n2036), .QN(n2031) );
  INVX0 U2042 ( .INP(n1964), .ZN(n2036) );
  XOR2X1 U2043 ( .IN1(n2037), .IN2(keyinput73), .Q(n1964) );
  OR2X1 U2044 ( .IN1(n2035), .IN2(n2034), .Q(n2037) );
  AO21X1 U2045 ( .IN1(n2038), .IN2(n2039), .IN3(n2040), .Q(n2035) );
  INVX0 U2046 ( .INP(n1962), .ZN(n2040) );
  XOR2X1 U2047 ( .IN1(n2041), .IN2(keyinput67), .Q(n1962) );
  OR2X1 U2048 ( .IN1(n2039), .IN2(n2038), .Q(n2041) );
  NAND2X0 U2049 ( .IN1(n1966), .IN2(n2042), .QN(n2039) );
  NAND3X0 U2050 ( .IN1(N409), .IN2(n2043), .IN3(N222), .QN(n2042) );
  AO21X1 U2051 ( .IN1(N222), .IN2(N409), .IN3(n2043), .Q(n1966) );
  NAND2X0 U2052 ( .IN1(n1967), .IN2(n2044), .QN(n2043) );
  NAND3X0 U2053 ( .IN1(n2045), .IN2(n2046), .IN3(n2047), .QN(n2044) );
  AO21X1 U2054 ( .IN1(n2045), .IN2(n2046), .IN3(n2047), .Q(n1967) );
  XNOR2X1 U2055 ( .IN1(n1973), .IN2(n1974), .Q(n2047) );
  NAND2X0 U2056 ( .IN1(N392), .IN2(N239), .QN(n1974) );
  XOR3X1 U2057 ( .IN1(keyinput51), .IN2(n2048), .IN3(n1971), .Q(n1973) );
  NAND2X0 U2058 ( .IN1(n2049), .IN2(n2050), .QN(n1971) );
  INVX0 U2059 ( .INP(n2051), .ZN(n2050) );
  AND2X1 U2060 ( .IN1(n2052), .IN2(n2053), .Q(n2038) );
  AO21X1 U2061 ( .IN1(n2054), .IN2(n2055), .IN3(n2056), .Q(n2052) );
  AND2X1 U2062 ( .IN1(N205), .IN2(N426), .Q(n2034) );
  INVX0 U2063 ( .INP(n2057), .ZN(n2032) );
  AND2X1 U2064 ( .IN1(N171), .IN2(N460), .Q(n2018) );
  XNOR2X1 U2065 ( .IN1(n2058), .IN2(keyinput13), .Q(n2005) );
  NAND2X0 U2066 ( .IN1(N137), .IN2(N494), .QN(n2058) );
  INVX0 U2067 ( .INP(n2059), .ZN(n2003) );
  NAND2X0 U2068 ( .IN1(n1982), .IN2(n2060), .QN(N6190) );
  NAND3X0 U2069 ( .IN1(n2061), .IN2(n2062), .IN3(n2063), .QN(n2060) );
  AO21X1 U2070 ( .IN1(n2061), .IN2(n2062), .IN3(n2063), .Q(n1982) );
  NAND2X0 U2071 ( .IN1(n1983), .IN2(n2064), .QN(n2063) );
  NAND3X0 U2072 ( .IN1(n2065), .IN2(n2066), .IN3(n2067), .QN(n2064) );
  AO21X1 U2073 ( .IN1(n2065), .IN2(n2066), .IN3(n2067), .Q(n1983) );
  XNOR2X1 U2074 ( .IN1(n1987), .IN2(n1988), .Q(n2067) );
  NAND2X0 U2075 ( .IN1(n2068), .IN2(n2069), .QN(n1988) );
  XNOR2X1 U2076 ( .IN1(n2070), .IN2(keyinput118), .Q(n2069) );
  NAND3X0 U2077 ( .IN1(n2071), .IN2(n1995), .IN3(n2072), .QN(n2070) );
  XNOR2X1 U2078 ( .IN1(keyinput119), .IN2(n2073), .Q(n2068) );
  AOI21X1 U2079 ( .IN1(n2074), .IN2(n2075), .IN3(n1989), .QN(n2073) );
  INVX0 U2080 ( .INP(n2072), .ZN(n1989) );
  NAND3X0 U2081 ( .IN1(n2071), .IN2(n1995), .IN3(n2076), .QN(n2072) );
  NAND2X0 U2082 ( .IN1(n2075), .IN2(n2074), .QN(n2076) );
  AO21X1 U2083 ( .IN1(N103), .IN2(N511), .IN3(n2077), .Q(n1995) );
  NAND3X0 U2084 ( .IN1(N511), .IN2(n2077), .IN3(N103), .QN(n2071) );
  NAND2X0 U2085 ( .IN1(n1996), .IN2(n2078), .QN(n2077) );
  NAND3X0 U2086 ( .IN1(n2079), .IN2(n2080), .IN3(n2081), .QN(n2078) );
  AO21X1 U2087 ( .IN1(n2079), .IN2(n2080), .IN3(n2081), .Q(n1996) );
  NAND2X0 U2088 ( .IN1(n2002), .IN2(n2082), .QN(n2081) );
  NAND3X0 U2089 ( .IN1(N494), .IN2(n2083), .IN3(N120), .QN(n2082) );
  AO21X1 U2090 ( .IN1(N120), .IN2(N494), .IN3(n2083), .Q(n2002) );
  AO21X1 U2091 ( .IN1(n2084), .IN2(n2085), .IN3(n2059), .Q(n2083) );
  NOR2X0 U2092 ( .IN1(n2085), .IN2(n2084), .QN(n2059) );
  NAND2X0 U2093 ( .IN1(n2009), .IN2(n2086), .QN(n2085) );
  NAND3X0 U2094 ( .IN1(N477), .IN2(n2087), .IN3(N137), .QN(n2086) );
  AO21X1 U2095 ( .IN1(N137), .IN2(N477), .IN3(n2087), .Q(n2009) );
  NAND2X0 U2096 ( .IN1(n2010), .IN2(n2088), .QN(n2087) );
  NAND3X0 U2097 ( .IN1(n2089), .IN2(n2090), .IN3(n2091), .QN(n2088) );
  AO21X1 U2098 ( .IN1(n2089), .IN2(n2090), .IN3(n2091), .Q(n2010) );
  NAND2X0 U2099 ( .IN1(n2015), .IN2(n2092), .QN(n2091) );
  NAND3X0 U2100 ( .IN1(N460), .IN2(n2093), .IN3(N154), .QN(n2092) );
  AO21X1 U2101 ( .IN1(N154), .IN2(N460), .IN3(n2093), .Q(n2015) );
  NAND2X0 U2102 ( .IN1(n2016), .IN2(n2094), .QN(n2093) );
  NAND3X0 U2103 ( .IN1(n2095), .IN2(n2096), .IN3(n2097), .QN(n2094) );
  AO21X1 U2104 ( .IN1(n2095), .IN2(n2096), .IN3(n2097), .Q(n2016) );
  NAND2X0 U2105 ( .IN1(n2022), .IN2(n2098), .QN(n2097) );
  NAND3X0 U2106 ( .IN1(N171), .IN2(N443), .IN3(n2099), .QN(n2098) );
  AO21X1 U2107 ( .IN1(N171), .IN2(N443), .IN3(n2099), .Q(n2022) );
  AOI21X1 U2108 ( .IN1(n2023), .IN2(n2100), .IN3(n2101), .QN(n2099) );
  XOR2X1 U2109 ( .IN1(n2102), .IN2(keyinput83), .Q(n2101) );
  NAND2X0 U2110 ( .IN1(n2103), .IN2(n2023), .QN(n2102) );
  INVX0 U2111 ( .INP(n2104), .ZN(n2103) );
  NAND2X0 U2112 ( .IN1(n2105), .IN2(n2106), .QN(n2100) );
  AO21X1 U2113 ( .IN1(n2105), .IN2(n2106), .IN3(n2104), .Q(n2023) );
  AO21X1 U2114 ( .IN1(n2107), .IN2(n2108), .IN3(n2033), .Q(n2104) );
  NOR2X0 U2115 ( .IN1(n2108), .IN2(n2107), .QN(n2033) );
  NAND2X0 U2116 ( .IN1(n2057), .IN2(n2109), .QN(n2108) );
  NAND3X0 U2117 ( .IN1(n2110), .IN2(n2111), .IN3(n2112), .QN(n2109) );
  AO21X1 U2118 ( .IN1(n2110), .IN2(n2111), .IN3(n2112), .Q(n2057) );
  NAND2X0 U2119 ( .IN1(n2053), .IN2(n2113), .QN(n2112) );
  NAND3X0 U2120 ( .IN1(N409), .IN2(n2114), .IN3(N205), .QN(n2113) );
  AO21X1 U2121 ( .IN1(N205), .IN2(N409), .IN3(n2114), .Q(n2053) );
  XNOR2X1 U2122 ( .IN1(n2056), .IN2(n2115), .Q(n2114) );
  AND2X1 U2123 ( .IN1(n2054), .IN2(n2055), .Q(n2115) );
  NAND2X0 U2124 ( .IN1(n2045), .IN2(n2116), .QN(n2056) );
  NAND3X0 U2125 ( .IN1(N222), .IN2(N392), .IN3(n2117), .QN(n2116) );
  AO21X1 U2126 ( .IN1(N222), .IN2(N392), .IN3(n2117), .Q(n2045) );
  XOR2X1 U2127 ( .IN1(n2118), .IN2(keyinput52), .Q(n2117) );
  NAND2X0 U2128 ( .IN1(n2046), .IN2(n2119), .QN(n2118) );
  NAND3X0 U2129 ( .IN1(n2120), .IN2(n2121), .IN3(n2122), .QN(n2119) );
  AO21X1 U2130 ( .IN1(n2120), .IN2(n2121), .IN3(n2122), .Q(n2046) );
  NAND3X0 U2131 ( .IN1(n2123), .IN2(n2049), .IN3(n2124), .QN(n2122) );
  NAND3X0 U2132 ( .IN1(n2048), .IN2(n2125), .IN3(n2126), .QN(n2124) );
  INVX0 U2133 ( .INP(n1972), .ZN(n2048) );
  NAND2X0 U2134 ( .IN1(N375), .IN2(N256), .QN(n1972) );
  AO221X1 U2135 ( .IN1(n2125), .IN2(n2127), .IN3(N375), .IN4(N239), .IN5(n2051), .Q(n2049) );
  NAND3X0 U2136 ( .IN1(N375), .IN2(N239), .IN3(n2051), .QN(n2123) );
  NOR2X0 U2137 ( .IN1(n2127), .IN2(n2125), .QN(n2051) );
  AOI21X1 U2138 ( .IN1(n2128), .IN2(n2129), .IN3(n2130), .QN(n2125) );
  NOR2X0 U2139 ( .IN1(n2131), .IN2(n1976), .QN(n2127) );
  INVX0 U2140 ( .INP(N256), .ZN(n1976) );
  XNOR2X1 U2141 ( .IN1(n2132), .IN2(keyinput16), .Q(n2107) );
  NAND2X0 U2142 ( .IN1(N188), .IN2(N426), .QN(n2132) );
  INVX0 U2143 ( .INP(n2133), .ZN(n2105) );
  XOR2X1 U2144 ( .IN1(n2134), .IN2(keyinput9), .Q(n1987) );
  NAND2X0 U2145 ( .IN1(N86), .IN2(N528), .QN(n2134) );
  INVX0 U2146 ( .INP(n2135), .ZN(n2062) );
  AO21X1 U2147 ( .IN1(n2136), .IN2(n2137), .IN3(n2135), .Q(N6180) );
  NOR2X0 U2148 ( .IN1(n2137), .IN2(n2136), .QN(n2135) );
  NAND2X0 U2149 ( .IN1(n2061), .IN2(n2138), .QN(n2137) );
  NAND3X0 U2150 ( .IN1(n2139), .IN2(n2140), .IN3(n2141), .QN(n2138) );
  AO21X1 U2151 ( .IN1(n2139), .IN2(n2140), .IN3(n2141), .Q(n2061) );
  NAND2X0 U2152 ( .IN1(n2065), .IN2(n2142), .QN(n2141) );
  NAND4X0 U2153 ( .IN1(N69), .IN2(N528), .IN3(n2143), .IN4(n2144), .QN(n2142)
         );
  AO22X1 U2154 ( .IN1(N69), .IN2(N528), .IN3(n2143), .IN4(n2144), .Q(n2065) );
  NAND2X0 U2155 ( .IN1(n2145), .IN2(n2066), .QN(n2144) );
  INVX0 U2156 ( .INP(n2146), .ZN(n2145) );
  XOR2X1 U2157 ( .IN1(keyinput120), .IN2(n2147), .Q(n2143) );
  OA21X1 U2158 ( .IN1(n2148), .IN2(n2149), .IN3(n2066), .Q(n2147) );
  AO21X1 U2159 ( .IN1(n2150), .IN2(n2151), .IN3(n2146), .Q(n2066) );
  NAND2X0 U2160 ( .IN1(n2152), .IN2(n2075), .QN(n2146) );
  AO21X1 U2161 ( .IN1(N86), .IN2(N511), .IN3(n2153), .Q(n2075) );
  NAND3X0 U2162 ( .IN1(N86), .IN2(N511), .IN3(n2153), .QN(n2152) );
  XOR2X1 U2163 ( .IN1(n2154), .IN2(keyinput112), .Q(n2153) );
  NAND2X0 U2164 ( .IN1(n2074), .IN2(n2155), .QN(n2154) );
  NAND3X0 U2165 ( .IN1(n2156), .IN2(n2157), .IN3(n2158), .QN(n2155) );
  AO21X1 U2166 ( .IN1(n2156), .IN2(n2157), .IN3(n2158), .Q(n2074) );
  NAND2X0 U2167 ( .IN1(n2079), .IN2(n2159), .QN(n2158) );
  NAND3X0 U2168 ( .IN1(N494), .IN2(n2160), .IN3(N103), .QN(n2159) );
  AO21X1 U2169 ( .IN1(N103), .IN2(N494), .IN3(n2160), .Q(n2079) );
  NAND2X0 U2170 ( .IN1(n2080), .IN2(n2161), .QN(n2160) );
  NAND3X0 U2171 ( .IN1(n2162), .IN2(n2163), .IN3(n2164), .QN(n2161) );
  AO21X1 U2172 ( .IN1(n2162), .IN2(n2163), .IN3(n2164), .Q(n2080) );
  OA21X1 U2173 ( .IN1(n2165), .IN2(n2166), .IN3(n2167), .Q(n2164) );
  NAND2X0 U2174 ( .IN1(n2084), .IN2(n2168), .QN(n2163) );
  AND2X1 U2175 ( .IN1(n2169), .IN2(n2170), .Q(n2084) );
  XOR2X1 U2176 ( .IN1(n2171), .IN2(keyinput99), .Q(n2162) );
  NAND2X0 U2177 ( .IN1(n2169), .IN2(n2172), .QN(n2171) );
  NAND3X0 U2178 ( .IN1(n2172), .IN2(n2170), .IN3(n2168), .QN(n2169) );
  NAND3X0 U2179 ( .IN1(n2173), .IN2(n2174), .IN3(n2175), .QN(n2168) );
  AO21X1 U2180 ( .IN1(n2173), .IN2(n2174), .IN3(n2175), .Q(n2170) );
  NAND2X0 U2181 ( .IN1(n2089), .IN2(n2176), .QN(n2175) );
  NAND3X0 U2182 ( .IN1(N460), .IN2(n2177), .IN3(N137), .QN(n2176) );
  AO21X1 U2183 ( .IN1(N137), .IN2(N460), .IN3(n2177), .Q(n2089) );
  NAND2X0 U2184 ( .IN1(n2090), .IN2(n2178), .QN(n2177) );
  NAND3X0 U2185 ( .IN1(n2179), .IN2(n2180), .IN3(n2181), .QN(n2178) );
  AO21X1 U2186 ( .IN1(n2179), .IN2(n2180), .IN3(n2181), .Q(n2090) );
  AOI21X1 U2187 ( .IN1(n2182), .IN2(n2183), .IN3(n2184), .QN(n2181) );
  INVX0 U2188 ( .INP(n2185), .ZN(n2184) );
  NAND2X0 U2189 ( .IN1(n2186), .IN2(n2095), .QN(n2180) );
  XOR2X1 U2190 ( .IN1(n2187), .IN2(keyinput90), .Q(n2179) );
  NAND2X0 U2191 ( .IN1(n2095), .IN2(n2188), .QN(n2187) );
  NAND2X0 U2192 ( .IN1(n2186), .IN2(n2188), .QN(n2095) );
  NAND2X0 U2193 ( .IN1(N154), .IN2(N443), .QN(n2188) );
  AND2X1 U2194 ( .IN1(n2189), .IN2(n2096), .Q(n2186) );
  AO221X1 U2195 ( .IN1(n2190), .IN2(n2191), .IN3(n2192), .IN4(n2193), .IN5(
        n2133), .Q(n2096) );
  NOR2X0 U2196 ( .IN1(n2191), .IN2(n2190), .QN(n2133) );
  NAND3X0 U2197 ( .IN1(n2192), .IN2(n2193), .IN3(n2194), .QN(n2189) );
  XNOR2X1 U2198 ( .IN1(n2191), .IN2(n2190), .Q(n2194) );
  AND2X1 U2199 ( .IN1(N171), .IN2(N426), .Q(n2190) );
  NAND2X0 U2200 ( .IN1(n2106), .IN2(n2195), .QN(n2191) );
  NAND3X0 U2201 ( .IN1(n2196), .IN2(n2197), .IN3(n2198), .QN(n2195) );
  AO21X1 U2202 ( .IN1(n2196), .IN2(n2197), .IN3(n2198), .Q(n2106) );
  NAND2X0 U2203 ( .IN1(n2110), .IN2(n2199), .QN(n2198) );
  NAND3X0 U2204 ( .IN1(N409), .IN2(n2200), .IN3(N188), .QN(n2199) );
  AO21X1 U2205 ( .IN1(N188), .IN2(N409), .IN3(n2200), .Q(n2110) );
  NAND2X0 U2206 ( .IN1(n2111), .IN2(n2201), .QN(n2200) );
  NAND3X0 U2207 ( .IN1(n2202), .IN2(n2203), .IN3(n2204), .QN(n2201) );
  AO21X1 U2208 ( .IN1(n2202), .IN2(n2203), .IN3(n2204), .Q(n2111) );
  NAND2X0 U2209 ( .IN1(n2054), .IN2(n2205), .QN(n2204) );
  NAND3X0 U2210 ( .IN1(N392), .IN2(n2206), .IN3(N205), .QN(n2205) );
  AO21X1 U2211 ( .IN1(N205), .IN2(N392), .IN3(n2206), .Q(n2054) );
  NAND2X0 U2212 ( .IN1(n2055), .IN2(n2207), .QN(n2206) );
  NAND3X0 U2213 ( .IN1(n2208), .IN2(n2209), .IN3(n2210), .QN(n2207) );
  AO21X1 U2214 ( .IN1(n2208), .IN2(n2209), .IN3(n2210), .Q(n2055) );
  NAND2X0 U2215 ( .IN1(n2120), .IN2(n2211), .QN(n2210) );
  NAND3X0 U2216 ( .IN1(N375), .IN2(n2212), .IN3(N222), .QN(n2211) );
  AO21X1 U2217 ( .IN1(N222), .IN2(N375), .IN3(n2212), .Q(n2120) );
  NAND2X0 U2218 ( .IN1(n2121), .IN2(n2213), .QN(n2212) );
  NAND3X0 U2219 ( .IN1(n2214), .IN2(n2215), .IN3(n2216), .QN(n2213) );
  AO21X1 U2220 ( .IN1(n2214), .IN2(n2215), .IN3(n2216), .Q(n2121) );
  AO21X1 U2221 ( .IN1(n2217), .IN2(n2126), .IN3(n2130), .Q(n2216) );
  XOR2X1 U2222 ( .IN1(n2218), .IN2(keyinput44), .Q(n2130) );
  OR2X1 U2223 ( .IN1(n2217), .IN2(n2126), .Q(n2218) );
  AND2X1 U2224 ( .IN1(N358), .IN2(N239), .Q(n2126) );
  XNOR2X1 U2225 ( .IN1(n2129), .IN2(n2128), .Q(n2217) );
  XNOR2X1 U2226 ( .IN1(keyinput40), .IN2(n2219), .Q(n2128) );
  OA21X1 U2227 ( .IN1(n2220), .IN2(n2221), .IN3(n2222), .Q(n2219) );
  NAND2X0 U2228 ( .IN1(N341), .IN2(N256), .QN(n2129) );
  NAND2X0 U2229 ( .IN1(N120), .IN2(N477), .QN(n2172) );
  INVX0 U2230 ( .INP(n2150), .ZN(n2149) );
  XNOR2X1 U2231 ( .IN1(keyinput125), .IN2(n2223), .Q(n2136) );
  AOI21X1 U2232 ( .IN1(n2224), .IN2(n2225), .IN3(n2226), .QN(n2223) );
  INVX0 U2233 ( .INP(n2227), .ZN(n2226) );
  XOR3X1 U2234 ( .IN1(keyinput126), .IN2(n2224), .IN3(n2225), .Q(N6170) );
  NAND2X0 U2235 ( .IN1(n2228), .IN2(n2229), .QN(n2225) );
  AND2X1 U2236 ( .IN1(n2227), .IN2(n2230), .Q(n2224) );
  NAND3X0 U2237 ( .IN1(n2231), .IN2(n2232), .IN3(n2233), .QN(n2230) );
  AO21X1 U2238 ( .IN1(n2231), .IN2(n2232), .IN3(n2233), .Q(n2227) );
  NAND2X0 U2239 ( .IN1(n2139), .IN2(n2234), .QN(n2233) );
  NAND3X0 U2240 ( .IN1(N528), .IN2(n2235), .IN3(N52), .QN(n2234) );
  AO21X1 U2241 ( .IN1(N52), .IN2(N528), .IN3(n2235), .Q(n2139) );
  NAND2X0 U2242 ( .IN1(n2140), .IN2(n2236), .QN(n2235) );
  NAND3X0 U2243 ( .IN1(n2237), .IN2(n2238), .IN3(n2239), .QN(n2236) );
  AO21X1 U2244 ( .IN1(n2237), .IN2(n2238), .IN3(n2239), .Q(n2140) );
  NAND2X0 U2245 ( .IN1(n2150), .IN2(n2240), .QN(n2239) );
  NAND3X0 U2246 ( .IN1(N69), .IN2(N511), .IN3(n2241), .QN(n2240) );
  AO21X1 U2247 ( .IN1(N69), .IN2(N511), .IN3(n2241), .Q(n2150) );
  AOI21X1 U2248 ( .IN1(n2151), .IN2(n2242), .IN3(n2243), .QN(n2241) );
  XOR2X1 U2249 ( .IN1(n2244), .IN2(keyinput111), .Q(n2243) );
  OR2X1 U2250 ( .IN1(n2245), .IN2(n2148), .Q(n2244) );
  INVX0 U2251 ( .INP(n2151), .ZN(n2148) );
  NAND2X0 U2252 ( .IN1(n2246), .IN2(n2247), .QN(n2242) );
  AO21X1 U2253 ( .IN1(n2246), .IN2(n2247), .IN3(n2245), .Q(n2151) );
  NAND2X0 U2254 ( .IN1(n2156), .IN2(n2248), .QN(n2245) );
  NAND3X0 U2255 ( .IN1(N494), .IN2(n2249), .IN3(N86), .QN(n2248) );
  AO21X1 U2256 ( .IN1(N86), .IN2(N494), .IN3(n2249), .Q(n2156) );
  NAND2X0 U2257 ( .IN1(n2157), .IN2(n2250), .QN(n2249) );
  NAND3X0 U2258 ( .IN1(n2251), .IN2(n2252), .IN3(n2253), .QN(n2250) );
  AO21X1 U2259 ( .IN1(n2251), .IN2(n2252), .IN3(n2253), .Q(n2157) );
  NAND2X0 U2260 ( .IN1(n2167), .IN2(n2254), .QN(n2253) );
  NAND3X0 U2261 ( .IN1(N477), .IN2(n2255), .IN3(N103), .QN(n2254) );
  AO21X1 U2262 ( .IN1(N103), .IN2(N477), .IN3(n2255), .Q(n2167) );
  XNOR2X1 U2263 ( .IN1(n2165), .IN2(n2166), .Q(n2255) );
  AND2X1 U2264 ( .IN1(n2256), .IN2(n2257), .Q(n2166) );
  NAND2X0 U2265 ( .IN1(n2173), .IN2(n2258), .QN(n2165) );
  NAND3X0 U2266 ( .IN1(N460), .IN2(n2259), .IN3(N120), .QN(n2258) );
  AO21X1 U2267 ( .IN1(N120), .IN2(N460), .IN3(n2259), .Q(n2173) );
  NAND2X0 U2268 ( .IN1(n2174), .IN2(n2260), .QN(n2259) );
  NAND3X0 U2269 ( .IN1(n2261), .IN2(n2262), .IN3(n2263), .QN(n2260) );
  AO21X1 U2270 ( .IN1(n2261), .IN2(n2262), .IN3(n2263), .Q(n2174) );
  OAI21X1 U2271 ( .IN1(n2264), .IN2(n2265), .IN3(n2185), .QN(n2263) );
  XOR2X1 U2272 ( .IN1(n2266), .IN2(keyinput89), .Q(n2185) );
  NAND2X0 U2273 ( .IN1(n2265), .IN2(n2264), .QN(n2266) );
  XOR2X1 U2274 ( .IN1(n2182), .IN2(n2183), .Q(n2265) );
  NAND2X0 U2275 ( .IN1(n2267), .IN2(n2268), .QN(n2183) );
  AO21X1 U2276 ( .IN1(N154), .IN2(N426), .IN3(n2269), .Q(n2268) );
  INVX0 U2277 ( .INP(n2192), .ZN(n2269) );
  XOR2X1 U2278 ( .IN1(n2270), .IN2(keyinput80), .Q(n2267) );
  NAND3X0 U2279 ( .IN1(n2271), .IN2(n2193), .IN3(n2192), .QN(n2270) );
  NAND3X0 U2280 ( .IN1(n2271), .IN2(n2193), .IN3(n2272), .QN(n2192) );
  NAND2X0 U2281 ( .IN1(N154), .IN2(N426), .QN(n2272) );
  AO21X1 U2282 ( .IN1(n2273), .IN2(n2274), .IN3(n2275), .Q(n2193) );
  NAND3X0 U2283 ( .IN1(n2273), .IN2(n2274), .IN3(n2275), .QN(n2271) );
  NAND2X0 U2284 ( .IN1(n2196), .IN2(n2276), .QN(n2275) );
  NAND3X0 U2285 ( .IN1(N409), .IN2(n2277), .IN3(N171), .QN(n2276) );
  AO21X1 U2286 ( .IN1(N171), .IN2(N409), .IN3(n2277), .Q(n2196) );
  NAND2X0 U2287 ( .IN1(n2197), .IN2(n2278), .QN(n2277) );
  NAND3X0 U2288 ( .IN1(n2279), .IN2(n2280), .IN3(n2281), .QN(n2278) );
  AO21X1 U2289 ( .IN1(n2279), .IN2(n2280), .IN3(n2281), .Q(n2197) );
  NAND2X0 U2290 ( .IN1(n2202), .IN2(n2282), .QN(n2281) );
  NAND3X0 U2291 ( .IN1(N188), .IN2(N392), .IN3(n2283), .QN(n2282) );
  AO21X1 U2292 ( .IN1(N188), .IN2(N392), .IN3(n2283), .Q(n2202) );
  XOR2X1 U2293 ( .IN1(n2284), .IN2(keyinput57), .Q(n2283) );
  NAND2X0 U2294 ( .IN1(n2203), .IN2(n2285), .QN(n2284) );
  AO221X1 U2295 ( .IN1(n2286), .IN2(n2208), .IN3(n2287), .IN4(n2288), .IN5(
        n2289), .Q(n2285) );
  NAND3X0 U2296 ( .IN1(n2286), .IN2(n2208), .IN3(n2290), .QN(n2203) );
  AO21X1 U2297 ( .IN1(n2287), .IN2(n2288), .IN3(n2289), .Q(n2290) );
  INVX0 U2298 ( .INP(n2291), .ZN(n2289) );
  AO21X1 U2299 ( .IN1(N205), .IN2(N375), .IN3(n2292), .Q(n2208) );
  NAND3X0 U2300 ( .IN1(N375), .IN2(n2292), .IN3(N205), .QN(n2286) );
  NAND2X0 U2301 ( .IN1(n2209), .IN2(n2293), .QN(n2292) );
  NAND3X0 U2302 ( .IN1(n2294), .IN2(n2295), .IN3(n2296), .QN(n2293) );
  AO21X1 U2303 ( .IN1(n2294), .IN2(n2295), .IN3(n2296), .Q(n2209) );
  NAND2X0 U2304 ( .IN1(n2214), .IN2(n2297), .QN(n2296) );
  NAND3X0 U2305 ( .IN1(N358), .IN2(n2298), .IN3(N222), .QN(n2297) );
  AO21X1 U2306 ( .IN1(N222), .IN2(N358), .IN3(n2298), .Q(n2214) );
  NAND2X0 U2307 ( .IN1(n2215), .IN2(n2299), .QN(n2298) );
  NAND3X0 U2308 ( .IN1(n2300), .IN2(n2301), .IN3(n2302), .QN(n2299) );
  AO21X1 U2309 ( .IN1(n2300), .IN2(n2301), .IN3(n2302), .Q(n2215) );
  XNOR2X1 U2310 ( .IN1(n2220), .IN2(n2221), .Q(n2302) );
  NAND2X0 U2311 ( .IN1(n2222), .IN2(n2303), .QN(n2221) );
  NAND4X0 U2312 ( .IN1(N324), .IN2(N256), .IN3(n2304), .IN4(n2305), .QN(n2303)
         );
  AO22X1 U2313 ( .IN1(n2306), .IN2(n2304), .IN3(N324), .IN4(N256), .Q(n2222)
         );
  AND2X1 U2314 ( .IN1(N341), .IN2(N239), .Q(n2220) );
  NAND2X0 U2315 ( .IN1(n2307), .IN2(n2308), .QN(n2182) );
  NAND2X0 U2316 ( .IN1(N137), .IN2(N443), .QN(n2264) );
  INVX0 U2317 ( .INP(n2309), .ZN(n2262) );
  XNOR2X1 U2318 ( .IN1(n2310), .IN2(keyinput124), .Q(N6160) );
  NAND2X0 U2319 ( .IN1(n2311), .IN2(n2229), .QN(n2310) );
  NAND3X0 U2320 ( .IN1(n2312), .IN2(n2228), .IN3(n2313), .QN(n2229) );
  NAND2X0 U2321 ( .IN1(n2314), .IN2(n2315), .QN(n2313) );
  NAND3X0 U2322 ( .IN1(n2316), .IN2(n2315), .IN3(n2314), .QN(n2311) );
  NAND2X0 U2323 ( .IN1(n2312), .IN2(n2228), .QN(n2316) );
  AO21X1 U2324 ( .IN1(n2317), .IN2(n2318), .IN3(n2319), .Q(n2228) );
  NAND3X0 U2325 ( .IN1(n2317), .IN2(n2318), .IN3(n2319), .QN(n2312) );
  NAND2X0 U2326 ( .IN1(n2231), .IN2(n2320), .QN(n2319) );
  NAND3X0 U2327 ( .IN1(N528), .IN2(n2321), .IN3(N35), .QN(n2320) );
  AO21X1 U2328 ( .IN1(N35), .IN2(N528), .IN3(n2321), .Q(n2231) );
  NAND2X0 U2329 ( .IN1(n2232), .IN2(n2322), .QN(n2321) );
  NAND3X0 U2330 ( .IN1(n2323), .IN2(n2324), .IN3(n2325), .QN(n2322) );
  AO21X1 U2331 ( .IN1(n2323), .IN2(n2324), .IN3(n2325), .Q(n2232) );
  NAND2X0 U2332 ( .IN1(n2237), .IN2(n2326), .QN(n2325) );
  NAND3X0 U2333 ( .IN1(N511), .IN2(n2327), .IN3(N52), .QN(n2326) );
  AO21X1 U2334 ( .IN1(N52), .IN2(N511), .IN3(n2327), .Q(n2237) );
  NAND2X0 U2335 ( .IN1(n2238), .IN2(n2328), .QN(n2327) );
  NAND3X0 U2336 ( .IN1(n2329), .IN2(n2330), .IN3(n2331), .QN(n2328) );
  AO21X1 U2337 ( .IN1(n2329), .IN2(n2330), .IN3(n2331), .Q(n2238) );
  NAND2X0 U2338 ( .IN1(n2246), .IN2(n2332), .QN(n2331) );
  NAND3X0 U2339 ( .IN1(N494), .IN2(n2333), .IN3(N69), .QN(n2332) );
  AO21X1 U2340 ( .IN1(N69), .IN2(N494), .IN3(n2333), .Q(n2246) );
  NAND2X0 U2341 ( .IN1(n2247), .IN2(n2334), .QN(n2333) );
  NAND3X0 U2342 ( .IN1(n2335), .IN2(n2336), .IN3(n2337), .QN(n2334) );
  AO21X1 U2343 ( .IN1(n2335), .IN2(n2336), .IN3(n2337), .Q(n2247) );
  NAND2X0 U2344 ( .IN1(n2251), .IN2(n2338), .QN(n2337) );
  NAND3X0 U2345 ( .IN1(N477), .IN2(n2339), .IN3(N86), .QN(n2338) );
  AO21X1 U2346 ( .IN1(N86), .IN2(N477), .IN3(n2339), .Q(n2251) );
  NAND2X0 U2347 ( .IN1(n2252), .IN2(n2340), .QN(n2339) );
  NAND3X0 U2348 ( .IN1(n2341), .IN2(n2342), .IN3(n2343), .QN(n2340) );
  AO21X1 U2349 ( .IN1(n2341), .IN2(n2342), .IN3(n2343), .Q(n2252) );
  NAND2X0 U2350 ( .IN1(n2257), .IN2(n2344), .QN(n2343) );
  NAND3X0 U2351 ( .IN1(N460), .IN2(n2345), .IN3(N103), .QN(n2344) );
  AO21X1 U2352 ( .IN1(N103), .IN2(N460), .IN3(n2345), .Q(n2257) );
  NAND2X0 U2353 ( .IN1(n2256), .IN2(n2346), .QN(n2345) );
  NAND3X0 U2354 ( .IN1(n2347), .IN2(n2348), .IN3(n2349), .QN(n2346) );
  AO21X1 U2355 ( .IN1(n2347), .IN2(n2348), .IN3(n2349), .Q(n2256) );
  AO21X1 U2356 ( .IN1(n2350), .IN2(n2351), .IN3(n2309), .Q(n2349) );
  NOR2X0 U2357 ( .IN1(n2351), .IN2(n2350), .QN(n2309) );
  XNOR2X1 U2358 ( .IN1(n2352), .IN2(keyinput11), .Q(n2351) );
  NAND2X0 U2359 ( .IN1(N120), .IN2(N443), .QN(n2352) );
  XNOR2X1 U2360 ( .IN1(keyinput88), .IN2(n2353), .Q(n2350) );
  AND2X1 U2361 ( .IN1(n2261), .IN2(n2354), .Q(n2353) );
  NAND3X0 U2362 ( .IN1(n2355), .IN2(n2356), .IN3(n2357), .QN(n2354) );
  AO21X1 U2363 ( .IN1(n2355), .IN2(n2356), .IN3(n2357), .Q(n2261) );
  NAND2X0 U2364 ( .IN1(n2308), .IN2(n2358), .QN(n2357) );
  NAND3X0 U2365 ( .IN1(N426), .IN2(n2359), .IN3(N137), .QN(n2358) );
  AO21X1 U2366 ( .IN1(N137), .IN2(N426), .IN3(n2359), .Q(n2308) );
  NAND2X0 U2367 ( .IN1(n2307), .IN2(n2360), .QN(n2359) );
  NAND3X0 U2368 ( .IN1(n2361), .IN2(n2362), .IN3(n2363), .QN(n2360) );
  AO21X1 U2369 ( .IN1(n2361), .IN2(n2362), .IN3(n2363), .Q(n2307) );
  NAND2X0 U2370 ( .IN1(n2273), .IN2(n2364), .QN(n2363) );
  NAND3X0 U2371 ( .IN1(N409), .IN2(n2365), .IN3(N154), .QN(n2364) );
  AO21X1 U2372 ( .IN1(N154), .IN2(N409), .IN3(n2365), .Q(n2273) );
  NAND2X0 U2373 ( .IN1(n2274), .IN2(n2366), .QN(n2365) );
  NAND3X0 U2374 ( .IN1(n2367), .IN2(n2368), .IN3(n2369), .QN(n2366) );
  AO21X1 U2375 ( .IN1(n2367), .IN2(n2368), .IN3(n2369), .Q(n2274) );
  NAND2X0 U2376 ( .IN1(n2279), .IN2(n2370), .QN(n2369) );
  NAND3X0 U2377 ( .IN1(N392), .IN2(n2371), .IN3(N171), .QN(n2370) );
  AO21X1 U2378 ( .IN1(N171), .IN2(N392), .IN3(n2371), .Q(n2279) );
  NAND2X0 U2379 ( .IN1(n2280), .IN2(n2372), .QN(n2371) );
  NAND3X0 U2380 ( .IN1(n2373), .IN2(n2374), .IN3(n2375), .QN(n2372) );
  AO21X1 U2381 ( .IN1(n2373), .IN2(n2374), .IN3(n2375), .Q(n2280) );
  XNOR2X1 U2382 ( .IN1(n2287), .IN2(n2288), .Q(n2375) );
  XNOR2X1 U2383 ( .IN1(n2376), .IN2(keyinput15), .Q(n2288) );
  NAND2X0 U2384 ( .IN1(N188), .IN2(N375), .QN(n2376) );
  AND2X1 U2385 ( .IN1(n2291), .IN2(n2377), .Q(n2287) );
  NAND3X0 U2386 ( .IN1(n2378), .IN2(n2379), .IN3(n2380), .QN(n2377) );
  AO21X1 U2387 ( .IN1(n2378), .IN2(n2379), .IN3(n2380), .Q(n2291) );
  NAND2X0 U2388 ( .IN1(n2294), .IN2(n2381), .QN(n2380) );
  NAND3X0 U2389 ( .IN1(n2382), .IN2(n2383), .IN3(n2384), .QN(n2381) );
  AO21X1 U2390 ( .IN1(n2382), .IN2(n2383), .IN3(n2384), .Q(n2294) );
  XNOR2X1 U2391 ( .IN1(n2385), .IN2(keyinput19), .Q(n2384) );
  NAND2X0 U2392 ( .IN1(N205), .IN2(N358), .QN(n2385) );
  OR2X1 U2393 ( .IN1(n2386), .IN2(n2387), .Q(n2383) );
  XOR2X1 U2394 ( .IN1(keyinput43), .IN2(n2388), .Q(n2382) );
  AOI21X1 U2395 ( .IN1(n2389), .IN2(n2390), .IN3(n2387), .QN(n2388) );
  INVX0 U2396 ( .INP(n2295), .ZN(n2387) );
  AO21X1 U2397 ( .IN1(n2390), .IN2(n2389), .IN3(n2386), .Q(n2295) );
  NAND2X0 U2398 ( .IN1(n2300), .IN2(n2391), .QN(n2386) );
  NAND3X0 U2399 ( .IN1(N341), .IN2(n2392), .IN3(N222), .QN(n2391) );
  AO21X1 U2400 ( .IN1(N222), .IN2(N341), .IN3(n2392), .Q(n2300) );
  NAND2X0 U2401 ( .IN1(n2301), .IN2(n2393), .QN(n2392) );
  NAND3X0 U2402 ( .IN1(n2394), .IN2(n2395), .IN3(n2396), .QN(n2393) );
  AO21X1 U2403 ( .IN1(n2394), .IN2(n2395), .IN3(n2396), .Q(n2301) );
  NAND2X0 U2404 ( .IN1(n2304), .IN2(n2397), .QN(n2396) );
  NAND3X0 U2405 ( .IN1(N239), .IN2(n2398), .IN3(N324), .QN(n2397) );
  AO21X1 U2406 ( .IN1(N324), .IN2(N239), .IN3(n2398), .Q(n2304) );
  NAND2X0 U2407 ( .IN1(n2399), .IN2(n2305), .QN(n2398) );
  OR2X1 U2408 ( .IN1(N307), .IN2(n2306), .Q(n2305) );
  MUX21X1 U2409 ( .IN1(n2306), .IN2(n2400), .S(N256), .Q(n2399) );
  NAND2X0 U2410 ( .IN1(n2306), .IN2(N307), .QN(n2400) );
  AND2X1 U2411 ( .IN1(n2401), .IN2(n2402), .Q(n2306) );
  AO21X1 U2412 ( .IN1(N290), .IN2(N256), .IN3(n2403), .Q(n2401) );
  XOR2X1 U2413 ( .IN1(n2314), .IN2(n2315), .Q(N6150) );
  NAND2X0 U2414 ( .IN1(n2317), .IN2(n2404), .QN(n2315) );
  NAND3X0 U2415 ( .IN1(N528), .IN2(n2405), .IN3(N18), .QN(n2404) );
  AO21X1 U2416 ( .IN1(N18), .IN2(N528), .IN3(n2405), .Q(n2317) );
  NAND2X0 U2417 ( .IN1(n2318), .IN2(n2406), .QN(n2405) );
  NAND3X0 U2418 ( .IN1(n2407), .IN2(n2408), .IN3(n2409), .QN(n2406) );
  AO21X1 U2419 ( .IN1(n2407), .IN2(n2408), .IN3(n2409), .Q(n2318) );
  NAND2X0 U2420 ( .IN1(n2323), .IN2(n2410), .QN(n2409) );
  NAND4X0 U2421 ( .IN1(n2411), .IN2(N35), .IN3(N511), .IN4(n2412), .QN(n2410)
         );
  AO22X1 U2422 ( .IN1(N35), .IN2(N511), .IN3(n2411), .IN4(n2412), .Q(n2323) );
  NAND2X0 U2423 ( .IN1(n2413), .IN2(n2324), .QN(n2412) );
  XOR2X1 U2424 ( .IN1(n2414), .IN2(keyinput116), .Q(n2411) );
  NAND2X0 U2425 ( .IN1(n2415), .IN2(n2324), .QN(n2414) );
  NAND2X0 U2426 ( .IN1(n2413), .IN2(n2415), .QN(n2324) );
  AND2X1 U2427 ( .IN1(n2329), .IN2(n2416), .Q(n2413) );
  NAND3X0 U2428 ( .IN1(N494), .IN2(n2417), .IN3(N52), .QN(n2416) );
  AO21X1 U2429 ( .IN1(N52), .IN2(N494), .IN3(n2417), .Q(n2329) );
  NAND2X0 U2430 ( .IN1(n2330), .IN2(n2418), .QN(n2417) );
  NAND3X0 U2431 ( .IN1(n2419), .IN2(n2420), .IN3(n2421), .QN(n2418) );
  AO21X1 U2432 ( .IN1(n2419), .IN2(n2420), .IN3(n2421), .Q(n2330) );
  XOR2X1 U2433 ( .IN1(n2422), .IN2(keyinput106), .Q(n2421) );
  NAND2X0 U2434 ( .IN1(n2335), .IN2(n2423), .QN(n2422) );
  NAND3X0 U2435 ( .IN1(N477), .IN2(n2424), .IN3(N69), .QN(n2423) );
  AO21X1 U2436 ( .IN1(N69), .IN2(N477), .IN3(n2424), .Q(n2335) );
  NAND2X0 U2437 ( .IN1(n2336), .IN2(n2425), .QN(n2424) );
  AO221X1 U2438 ( .IN1(n2426), .IN2(n2341), .IN3(n2427), .IN4(n2428), .IN5(
        n2429), .Q(n2425) );
  NAND3X0 U2439 ( .IN1(n2426), .IN2(n2341), .IN3(n2430), .QN(n2336) );
  AO21X1 U2440 ( .IN1(n2427), .IN2(n2428), .IN3(n2429), .Q(n2430) );
  INVX0 U2441 ( .INP(n2431), .ZN(n2429) );
  AO21X1 U2442 ( .IN1(N86), .IN2(N460), .IN3(n2432), .Q(n2341) );
  NAND3X0 U2443 ( .IN1(N460), .IN2(n2432), .IN3(N86), .QN(n2426) );
  NAND2X0 U2444 ( .IN1(n2342), .IN2(n2433), .QN(n2432) );
  NAND3X0 U2445 ( .IN1(n2434), .IN2(n2435), .IN3(n2436), .QN(n2433) );
  AO21X1 U2446 ( .IN1(n2434), .IN2(n2435), .IN3(n2436), .Q(n2342) );
  NAND2X0 U2447 ( .IN1(n2347), .IN2(n2437), .QN(n2436) );
  NAND3X0 U2448 ( .IN1(N103), .IN2(N443), .IN3(n2438), .QN(n2437) );
  AO21X1 U2449 ( .IN1(N103), .IN2(N443), .IN3(n2438), .Q(n2347) );
  AND2X1 U2450 ( .IN1(n2439), .IN2(n2440), .Q(n2438) );
  AO21X1 U2451 ( .IN1(n2441), .IN2(n2442), .IN3(n2443), .Q(n2440) );
  XOR2X1 U2452 ( .IN1(keyinput87), .IN2(n2444), .Q(n2439) );
  NOR2X0 U2453 ( .IN1(n2443), .IN2(n2445), .QN(n2444) );
  INVX0 U2454 ( .INP(n2348), .ZN(n2443) );
  AO21X1 U2455 ( .IN1(n2441), .IN2(n2442), .IN3(n2445), .Q(n2348) );
  NAND2X0 U2456 ( .IN1(n2446), .IN2(n2355), .QN(n2445) );
  AO21X1 U2457 ( .IN1(N120), .IN2(N426), .IN3(n2447), .Q(n2355) );
  NAND3X0 U2458 ( .IN1(N426), .IN2(n2447), .IN3(N120), .QN(n2446) );
  XNOR2X1 U2459 ( .IN1(keyinput79), .IN2(n2448), .Q(n2447) );
  AO21X1 U2460 ( .IN1(n2449), .IN2(n2356), .IN3(n2450), .Q(n2448) );
  XOR2X1 U2461 ( .IN1(keyinput77), .IN2(n2451), .Q(n2450) );
  NOR2X0 U2462 ( .IN1(n2452), .IN2(n2453), .QN(n2451) );
  INVX0 U2463 ( .INP(n2356), .ZN(n2453) );
  OA21X1 U2464 ( .IN1(n2454), .IN2(n2455), .IN3(n2456), .Q(n2452) );
  AO21X1 U2465 ( .IN1(n2456), .IN2(n2457), .IN3(n2458), .Q(n2356) );
  OR2X1 U2466 ( .IN1(n2455), .IN2(n2454), .Q(n2457) );
  INVX0 U2467 ( .INP(n2458), .ZN(n2449) );
  NAND2X0 U2468 ( .IN1(n2361), .IN2(n2459), .QN(n2458) );
  NAND3X0 U2469 ( .IN1(N137), .IN2(N409), .IN3(n2460), .QN(n2459) );
  AO21X1 U2470 ( .IN1(N137), .IN2(N409), .IN3(n2460), .Q(n2361) );
  AND2X1 U2471 ( .IN1(n2461), .IN2(n2462), .Q(n2460) );
  AO21X1 U2472 ( .IN1(n2463), .IN2(n2464), .IN3(n2465), .Q(n2462) );
  XOR2X1 U2473 ( .IN1(n2466), .IN2(keyinput66), .Q(n2461) );
  OR2X1 U2474 ( .IN1(n2467), .IN2(n2465), .Q(n2466) );
  INVX0 U2475 ( .INP(n2362), .ZN(n2465) );
  AO21X1 U2476 ( .IN1(n2463), .IN2(n2464), .IN3(n2467), .Q(n2362) );
  INVX0 U2477 ( .INP(n2468), .ZN(n2464) );
  NAND2X0 U2478 ( .IN1(n2469), .IN2(n2367), .QN(n2467) );
  NAND3X0 U2479 ( .IN1(n2470), .IN2(n2368), .IN3(n2471), .QN(n2367) );
  NAND2X0 U2480 ( .IN1(N154), .IN2(N392), .QN(n2471) );
  NAND3X0 U2481 ( .IN1(N392), .IN2(n2472), .IN3(N154), .QN(n2469) );
  NAND2X0 U2482 ( .IN1(n2470), .IN2(n2368), .QN(n2472) );
  AO21X1 U2483 ( .IN1(n2473), .IN2(n2474), .IN3(n2475), .Q(n2368) );
  NAND3X0 U2484 ( .IN1(n2473), .IN2(n2474), .IN3(n2475), .QN(n2470) );
  NAND2X0 U2485 ( .IN1(n2373), .IN2(n2476), .QN(n2475) );
  NAND3X0 U2486 ( .IN1(N375), .IN2(n2477), .IN3(N171), .QN(n2476) );
  AO21X1 U2487 ( .IN1(N171), .IN2(N375), .IN3(n2477), .Q(n2373) );
  NAND2X0 U2488 ( .IN1(n2374), .IN2(n2478), .QN(n2477) );
  NAND3X0 U2489 ( .IN1(n2479), .IN2(n2480), .IN3(n2481), .QN(n2478) );
  AO21X1 U2490 ( .IN1(n2479), .IN2(n2480), .IN3(n2481), .Q(n2374) );
  NAND2X0 U2491 ( .IN1(n2378), .IN2(n2482), .QN(n2481) );
  NAND3X0 U2492 ( .IN1(N358), .IN2(n2483), .IN3(N188), .QN(n2482) );
  AO21X1 U2493 ( .IN1(N188), .IN2(N358), .IN3(n2483), .Q(n2378) );
  NAND2X0 U2494 ( .IN1(n2379), .IN2(n2484), .QN(n2483) );
  NAND3X0 U2495 ( .IN1(n2485), .IN2(n2486), .IN3(n2487), .QN(n2484) );
  AO21X1 U2496 ( .IN1(n2485), .IN2(n2486), .IN3(n2487), .Q(n2379) );
  AND2X1 U2497 ( .IN1(n2488), .IN2(n2489), .Q(n2487) );
  AO21X1 U2498 ( .IN1(n2490), .IN2(n2491), .IN3(n2492), .Q(n2488) );
  NAND2X0 U2499 ( .IN1(n2493), .IN2(n2390), .QN(n2486) );
  XNOR2X1 U2500 ( .IN1(n2494), .IN2(keyinput42), .Q(n2485) );
  NAND2X0 U2501 ( .IN1(n2390), .IN2(n2495), .QN(n2494) );
  NAND2X0 U2502 ( .IN1(n2493), .IN2(n2495), .QN(n2390) );
  NAND2X0 U2503 ( .IN1(N205), .IN2(N341), .QN(n2495) );
  AND2X1 U2504 ( .IN1(n2389), .IN2(n2496), .Q(n2493) );
  NAND3X0 U2505 ( .IN1(n2497), .IN2(n2498), .IN3(n2499), .QN(n2496) );
  AO21X1 U2506 ( .IN1(n2497), .IN2(n2498), .IN3(n2499), .Q(n2389) );
  NAND2X0 U2507 ( .IN1(n2394), .IN2(n2500), .QN(n2499) );
  NAND3X0 U2508 ( .IN1(N324), .IN2(n2501), .IN3(N222), .QN(n2500) );
  AO21X1 U2509 ( .IN1(N222), .IN2(N324), .IN3(n2501), .Q(n2394) );
  NAND2X0 U2510 ( .IN1(n2395), .IN2(n2502), .QN(n2501) );
  NAND3X0 U2511 ( .IN1(n2503), .IN2(n2504), .IN3(n2505), .QN(n2502) );
  AO21X1 U2512 ( .IN1(n2503), .IN2(n2504), .IN3(n2505), .Q(n2395) );
  NAND2X0 U2513 ( .IN1(n2402), .IN2(n2506), .QN(n2505) );
  NAND3X0 U2514 ( .IN1(N307), .IN2(N239), .IN3(n2507), .QN(n2506) );
  AO21X1 U2515 ( .IN1(N307), .IN2(N239), .IN3(n2507), .Q(n2402) );
  XOR2X1 U2516 ( .IN1(n2508), .IN2(n2403), .Q(n2507) );
  AND3X1 U2517 ( .IN1(N239), .IN2(n2509), .IN3(N290), .Q(n2403) );
  NAND2X0 U2518 ( .IN1(N290), .IN2(N256), .QN(n2508) );
  INVX0 U2519 ( .INP(n2510), .ZN(n2504) );
  AO22X1 U2520 ( .IN1(n2511), .IN2(n2512), .IN3(n2513), .IN4(n2514), .Q(n2415)
         );
  OA21X1 U2521 ( .IN1(n2515), .IN2(n2516), .IN3(n2517), .Q(n2314) );
  AND2X1 U2522 ( .IN1(N1), .IN2(N528), .Q(n2516) );
  XOR2X1 U2523 ( .IN1(n2515), .IN2(n2518), .Q(N6123) );
  NAND2X0 U2524 ( .IN1(N1), .IN2(N528), .QN(n2518) );
  NAND2X0 U2525 ( .IN1(n2517), .IN2(n2519), .QN(n2515) );
  NAND3X0 U2526 ( .IN1(n2520), .IN2(n2521), .IN3(n2522), .QN(n2519) );
  AO21X1 U2527 ( .IN1(n2520), .IN2(n2521), .IN3(n2522), .Q(n2517) );
  NAND2X0 U2528 ( .IN1(n2407), .IN2(n2523), .QN(n2522) );
  NAND3X0 U2529 ( .IN1(N511), .IN2(n2524), .IN3(N18), .QN(n2523) );
  AO21X1 U2530 ( .IN1(N18), .IN2(N511), .IN3(n2524), .Q(n2407) );
  NAND2X0 U2531 ( .IN1(n2408), .IN2(n2525), .QN(n2524) );
  NAND3X0 U2532 ( .IN1(n2526), .IN2(n2527), .IN3(n2528), .QN(n2525) );
  AO21X1 U2533 ( .IN1(n2526), .IN2(n2527), .IN3(n2528), .Q(n2408) );
  XNOR2X1 U2534 ( .IN1(n2513), .IN2(n2514), .Q(n2528) );
  NAND2X0 U2535 ( .IN1(N35), .IN2(N494), .QN(n2514) );
  XOR2X1 U2536 ( .IN1(n2511), .IN2(n2512), .Q(n2513) );
  XOR2X1 U2537 ( .IN1(keyinput105), .IN2(n2529), .Q(n2512) );
  OA21X1 U2538 ( .IN1(n2530), .IN2(n2531), .IN3(n2532), .Q(n2529) );
  AND2X1 U2539 ( .IN1(n2419), .IN2(n2533), .Q(n2511) );
  NAND3X0 U2540 ( .IN1(N477), .IN2(n2534), .IN3(N52), .QN(n2533) );
  AO21X1 U2541 ( .IN1(N52), .IN2(N477), .IN3(n2534), .Q(n2419) );
  NAND2X0 U2542 ( .IN1(n2420), .IN2(n2535), .QN(n2534) );
  NAND3X0 U2543 ( .IN1(n2536), .IN2(n2537), .IN3(n2538), .QN(n2535) );
  AO21X1 U2544 ( .IN1(n2536), .IN2(n2537), .IN3(n2538), .Q(n2420) );
  XNOR2X1 U2545 ( .IN1(n2427), .IN2(n2428), .Q(n2538) );
  XOR2X1 U2546 ( .IN1(n2539), .IN2(keyinput8), .Q(n2428) );
  NAND2X0 U2547 ( .IN1(N69), .IN2(N460), .QN(n2539) );
  AND2X1 U2548 ( .IN1(n2431), .IN2(n2540), .Q(n2427) );
  NAND3X0 U2549 ( .IN1(n2541), .IN2(n2542), .IN3(n2543), .QN(n2540) );
  AO21X1 U2550 ( .IN1(n2541), .IN2(n2542), .IN3(n2543), .Q(n2431) );
  NAND2X0 U2551 ( .IN1(n2434), .IN2(n2544), .QN(n2543) );
  NAND3X0 U2552 ( .IN1(N443), .IN2(n2545), .IN3(N86), .QN(n2544) );
  AO21X1 U2553 ( .IN1(N86), .IN2(N443), .IN3(n2545), .Q(n2434) );
  NAND2X0 U2554 ( .IN1(n2435), .IN2(n2546), .QN(n2545) );
  NAND3X0 U2555 ( .IN1(n2547), .IN2(n2548), .IN3(n2549), .QN(n2546) );
  AO21X1 U2556 ( .IN1(n2547), .IN2(n2548), .IN3(n2549), .Q(n2435) );
  XOR2X1 U2557 ( .IN1(n2550), .IN2(keyinput86), .Q(n2549) );
  NAND2X0 U2558 ( .IN1(n2441), .IN2(n2551), .QN(n2550) );
  NAND3X0 U2559 ( .IN1(N426), .IN2(n2552), .IN3(N103), .QN(n2551) );
  AO21X1 U2560 ( .IN1(N103), .IN2(N426), .IN3(n2552), .Q(n2441) );
  NAND2X0 U2561 ( .IN1(n2442), .IN2(n2553), .QN(n2552) );
  NAND3X0 U2562 ( .IN1(n2554), .IN2(n2555), .IN3(n2556), .QN(n2553) );
  AO21X1 U2563 ( .IN1(n2554), .IN2(n2555), .IN3(n2556), .Q(n2442) );
  XOR3X1 U2564 ( .IN1(keyinput76), .IN2(n2454), .IN3(n2455), .Q(n2556) );
  NAND2X0 U2565 ( .IN1(n2456), .IN2(n2557), .QN(n2455) );
  NAND3X0 U2566 ( .IN1(n2558), .IN2(n2559), .IN3(n2560), .QN(n2557) );
  AO21X1 U2567 ( .IN1(n2558), .IN2(n2559), .IN3(n2560), .Q(n2456) );
  NAND2X0 U2568 ( .IN1(n2463), .IN2(n2561), .QN(n2560) );
  NAND3X0 U2569 ( .IN1(N392), .IN2(n2562), .IN3(N137), .QN(n2561) );
  AO21X1 U2570 ( .IN1(N137), .IN2(N392), .IN3(n2562), .Q(n2463) );
  AO21X1 U2571 ( .IN1(n2563), .IN2(n2564), .IN3(n2468), .Q(n2562) );
  NOR2X0 U2572 ( .IN1(n2564), .IN2(n2563), .QN(n2468) );
  NAND2X0 U2573 ( .IN1(n2473), .IN2(n2565), .QN(n2564) );
  NAND3X0 U2574 ( .IN1(N375), .IN2(n2566), .IN3(N154), .QN(n2565) );
  AO21X1 U2575 ( .IN1(N154), .IN2(N375), .IN3(n2566), .Q(n2473) );
  NAND2X0 U2576 ( .IN1(n2474), .IN2(n2567), .QN(n2566) );
  NAND3X0 U2577 ( .IN1(n2568), .IN2(n2569), .IN3(n2570), .QN(n2567) );
  AO21X1 U2578 ( .IN1(n2570), .IN2(n2569), .IN3(n2568), .Q(n2474) );
  NAND2X0 U2579 ( .IN1(n2479), .IN2(n2571), .QN(n2568) );
  NAND3X0 U2580 ( .IN1(N358), .IN2(n2572), .IN3(N171), .QN(n2571) );
  AO21X1 U2581 ( .IN1(N171), .IN2(N358), .IN3(n2572), .Q(n2479) );
  NAND2X0 U2582 ( .IN1(n2480), .IN2(n2573), .QN(n2572) );
  NAND3X0 U2583 ( .IN1(n2574), .IN2(n2575), .IN3(n2576), .QN(n2573) );
  AO21X1 U2584 ( .IN1(n2574), .IN2(n2575), .IN3(n2576), .Q(n2480) );
  NAND2X0 U2585 ( .IN1(n2489), .IN2(n2577), .QN(n2576) );
  NAND3X0 U2586 ( .IN1(N341), .IN2(n2578), .IN3(N188), .QN(n2577) );
  AO21X1 U2587 ( .IN1(N188), .IN2(N341), .IN3(n2578), .Q(n2489) );
  XOR2X1 U2588 ( .IN1(n2579), .IN2(n2492), .Q(n2578) );
  NAND2X0 U2589 ( .IN1(n2497), .IN2(n2580), .QN(n2492) );
  NAND3X0 U2590 ( .IN1(N324), .IN2(n2581), .IN3(N205), .QN(n2580) );
  AO21X1 U2591 ( .IN1(N205), .IN2(N324), .IN3(n2581), .Q(n2497) );
  NAND2X0 U2592 ( .IN1(n2498), .IN2(n2582), .QN(n2581) );
  NAND3X0 U2593 ( .IN1(n2583), .IN2(n2584), .IN3(n2585), .QN(n2582) );
  AO21X1 U2594 ( .IN1(n2583), .IN2(n2584), .IN3(n2585), .Q(n2498) );
  NAND2X0 U2595 ( .IN1(n2503), .IN2(n2586), .QN(n2585) );
  NAND3X0 U2596 ( .IN1(N307), .IN2(n2587), .IN3(N222), .QN(n2586) );
  AO21X1 U2597 ( .IN1(N222), .IN2(N307), .IN3(n2587), .Q(n2503) );
  AO21X1 U2598 ( .IN1(n2588), .IN2(n2589), .IN3(n2510), .Q(n2587) );
  NOR2X0 U2599 ( .IN1(n2589), .IN2(n2588), .QN(n2510) );
  XOR2X1 U2600 ( .IN1(n2509), .IN2(n2590), .Q(n2589) );
  AND2X1 U2601 ( .IN1(N239), .IN2(N290), .Q(n2590) );
  XNOR2X1 U2602 ( .IN1(n2591), .IN2(keyinput21), .Q(n2509) );
  NAND2X0 U2603 ( .IN1(N273), .IN2(N256), .QN(n2591) );
  INVX0 U2604 ( .INP(n2592), .ZN(n2588) );
  NAND2X0 U2605 ( .IN1(n2490), .IN2(n2491), .QN(n2579) );
  INVX0 U2606 ( .INP(n2593), .ZN(n2491) );
  AND2X1 U2607 ( .IN1(N120), .IN2(N409), .Q(n2454) );
  OA21X1 U2608 ( .IN1(n2594), .IN2(n2595), .IN3(n2596), .Q(N5971) );
  XOR2X1 U2609 ( .IN1(n2597), .IN2(keyinput122), .Q(n2596) );
  NAND2X0 U2610 ( .IN1(n2598), .IN2(n2521), .QN(n2597) );
  INVX0 U2611 ( .INP(n2594), .ZN(n2521) );
  XNOR2X1 U2612 ( .IN1(keyinput117), .IN2(n2599), .Q(n2598) );
  NOR2X0 U2613 ( .IN1(n2600), .IN2(n2595), .QN(n2594) );
  NOR2X0 U2614 ( .IN1(n2601), .IN2(n1908), .QN(n2595) );
  INVX0 U2615 ( .INP(N511), .ZN(n1908) );
  XOR2X1 U2616 ( .IN1(keyinput117), .IN2(n2599), .Q(n2600) );
  NAND2X0 U2617 ( .IN1(n2520), .IN2(n2602), .QN(n2599) );
  NAND3X0 U2618 ( .IN1(n2603), .IN2(n2604), .IN3(n2605), .QN(n2602) );
  AO21X1 U2619 ( .IN1(n2603), .IN2(n2604), .IN3(n2605), .Q(n2520) );
  NAND2X0 U2620 ( .IN1(n2526), .IN2(n2606), .QN(n2605) );
  NAND3X0 U2621 ( .IN1(N494), .IN2(n2607), .IN3(N18), .QN(n2606) );
  AO21X1 U2622 ( .IN1(N18), .IN2(N494), .IN3(n2607), .Q(n2526) );
  NAND2X0 U2623 ( .IN1(n2527), .IN2(n2608), .QN(n2607) );
  NAND3X0 U2624 ( .IN1(n2609), .IN2(n2610), .IN3(n2611), .QN(n2608) );
  AO21X1 U2625 ( .IN1(n2609), .IN2(n2610), .IN3(n2611), .Q(n2527) );
  XNOR2X1 U2626 ( .IN1(n2531), .IN2(n2530), .Q(n2611) );
  AND2X1 U2627 ( .IN1(N35), .IN2(N477), .Q(n2530) );
  NAND2X0 U2628 ( .IN1(n2532), .IN2(n2612), .QN(n2531) );
  NAND3X0 U2629 ( .IN1(n2613), .IN2(n2614), .IN3(n2615), .QN(n2612) );
  XOR2X1 U2630 ( .IN1(keyinput98), .IN2(n2616), .Q(n2532) );
  AOI21X1 U2631 ( .IN1(n2614), .IN2(n2613), .IN3(n2615), .QN(n2616) );
  NAND2X0 U2632 ( .IN1(n2536), .IN2(n2617), .QN(n2615) );
  NAND3X0 U2633 ( .IN1(N460), .IN2(n2618), .IN3(N52), .QN(n2617) );
  AO21X1 U2634 ( .IN1(N52), .IN2(N460), .IN3(n2618), .Q(n2536) );
  NAND2X0 U2635 ( .IN1(n2537), .IN2(n2619), .QN(n2618) );
  NAND3X0 U2636 ( .IN1(n2620), .IN2(n2621), .IN3(n2622), .QN(n2619) );
  AO21X1 U2637 ( .IN1(n2620), .IN2(n2621), .IN3(n2622), .Q(n2537) );
  NAND2X0 U2638 ( .IN1(n2541), .IN2(n2623), .QN(n2622) );
  NAND3X0 U2639 ( .IN1(N443), .IN2(n2624), .IN3(N69), .QN(n2623) );
  AO21X1 U2640 ( .IN1(N69), .IN2(N443), .IN3(n2624), .Q(n2541) );
  NAND2X0 U2641 ( .IN1(n2542), .IN2(n2625), .QN(n2624) );
  NAND3X0 U2642 ( .IN1(n2626), .IN2(n2627), .IN3(n2628), .QN(n2625) );
  AO21X1 U2643 ( .IN1(n2626), .IN2(n2627), .IN3(n2628), .Q(n2542) );
  NAND2X0 U2644 ( .IN1(n2547), .IN2(n2629), .QN(n2628) );
  NAND3X0 U2645 ( .IN1(N426), .IN2(n2630), .IN3(N86), .QN(n2629) );
  AO21X1 U2646 ( .IN1(N86), .IN2(N426), .IN3(n2630), .Q(n2547) );
  NAND2X0 U2647 ( .IN1(n2548), .IN2(n2631), .QN(n2630) );
  NAND3X0 U2648 ( .IN1(n2632), .IN2(n2633), .IN3(n2634), .QN(n2631) );
  AO21X1 U2649 ( .IN1(n2632), .IN2(n2633), .IN3(n2634), .Q(n2548) );
  OAI21X1 U2650 ( .IN1(n2635), .IN2(n2636), .IN3(n2554), .QN(n2634) );
  XOR2X1 U2651 ( .IN1(n2637), .IN2(keyinput72), .Q(n2554) );
  NAND2X0 U2652 ( .IN1(n2636), .IN2(n2635), .QN(n2637) );
  AO21X1 U2653 ( .IN1(n2638), .IN2(n2555), .IN3(n2639), .Q(n2636) );
  XNOR2X1 U2654 ( .IN1(keyinput69), .IN2(n2640), .Q(n2639) );
  AOI21X1 U2655 ( .IN1(n2641), .IN2(n2642), .IN3(n2643), .QN(n2640) );
  INVX0 U2656 ( .INP(n2555), .ZN(n2643) );
  AO21X1 U2657 ( .IN1(n2642), .IN2(n2641), .IN3(n2644), .Q(n2555) );
  XOR2X1 U2658 ( .IN1(n2645), .IN2(keyinput64), .Q(n2644) );
  XNOR2X1 U2659 ( .IN1(keyinput64), .IN2(n2645), .Q(n2638) );
  NAND2X0 U2660 ( .IN1(n2558), .IN2(n2646), .QN(n2645) );
  NAND3X0 U2661 ( .IN1(N392), .IN2(n2647), .IN3(N120), .QN(n2646) );
  AO21X1 U2662 ( .IN1(N120), .IN2(N392), .IN3(n2647), .Q(n2558) );
  OAI21X1 U2663 ( .IN1(n2648), .IN2(n2649), .IN3(n2559), .QN(n2647) );
  NAND2X0 U2664 ( .IN1(n2649), .IN2(n2648), .QN(n2559) );
  XNOR2X1 U2665 ( .IN1(keyinput55), .IN2(n2650), .Q(n2649) );
  OA21X1 U2666 ( .IN1(n2651), .IN2(n2652), .IN3(n2653), .Q(n2650) );
  NAND2X0 U2667 ( .IN1(n2654), .IN2(n2655), .QN(n2648) );
  AO21X1 U2668 ( .IN1(N137), .IN2(N375), .IN3(n2656), .Q(n2655) );
  INVX0 U2669 ( .INP(n2657), .ZN(n2656) );
  XOR2X1 U2670 ( .IN1(n2658), .IN2(keyinput56), .Q(n2654) );
  NAND2X0 U2671 ( .IN1(n2563), .IN2(n2659), .QN(n2658) );
  AND2X1 U2672 ( .IN1(n2657), .IN2(n2660), .Q(n2563) );
  NAND3X0 U2673 ( .IN1(n2659), .IN2(n2660), .IN3(n2661), .QN(n2657) );
  NAND2X0 U2674 ( .IN1(N137), .IN2(N375), .QN(n2661) );
  AO21X1 U2675 ( .IN1(n2662), .IN2(n2663), .IN3(n2664), .Q(n2660) );
  NAND3X0 U2676 ( .IN1(n2662), .IN2(n2663), .IN3(n2664), .QN(n2659) );
  NAND2X0 U2677 ( .IN1(n2570), .IN2(n2665), .QN(n2664) );
  NAND3X0 U2678 ( .IN1(N358), .IN2(n2666), .IN3(N154), .QN(n2665) );
  XNOR2X1 U2679 ( .IN1(keyinput47), .IN2(n2667), .Q(n2570) );
  AOI21X1 U2680 ( .IN1(N358), .IN2(N154), .IN3(n2666), .QN(n2667) );
  NAND2X0 U2681 ( .IN1(n2569), .IN2(n2668), .QN(n2666) );
  NAND3X0 U2682 ( .IN1(n2669), .IN2(n2670), .IN3(n2671), .QN(n2668) );
  AO21X1 U2683 ( .IN1(n2669), .IN2(n2670), .IN3(n2671), .Q(n2569) );
  NAND2X0 U2684 ( .IN1(n2574), .IN2(n2672), .QN(n2671) );
  NAND3X0 U2685 ( .IN1(N341), .IN2(n2673), .IN3(N171), .QN(n2672) );
  AO21X1 U2686 ( .IN1(N171), .IN2(N341), .IN3(n2673), .Q(n2574) );
  NAND2X0 U2687 ( .IN1(n2575), .IN2(n2674), .QN(n2673) );
  NAND3X0 U2688 ( .IN1(n2675), .IN2(n2676), .IN3(n2677), .QN(n2674) );
  AO21X1 U2689 ( .IN1(n2675), .IN2(n2676), .IN3(n2677), .Q(n2575) );
  NAND2X0 U2690 ( .IN1(n2490), .IN2(n2678), .QN(n2677) );
  NAND3X0 U2691 ( .IN1(N324), .IN2(n2679), .IN3(N188), .QN(n2678) );
  AO21X1 U2692 ( .IN1(N188), .IN2(N324), .IN3(n2679), .Q(n2490) );
  AO21X1 U2693 ( .IN1(n2680), .IN2(n2681), .IN3(n2593), .Q(n2679) );
  NOR2X0 U2694 ( .IN1(n2681), .IN2(n2680), .QN(n2593) );
  NAND2X0 U2695 ( .IN1(n2583), .IN2(n2682), .QN(n2681) );
  NAND3X0 U2696 ( .IN1(N307), .IN2(n2683), .IN3(N205), .QN(n2682) );
  AO21X1 U2697 ( .IN1(N205), .IN2(N307), .IN3(n2683), .Q(n2583) );
  AO21X1 U2698 ( .IN1(n2684), .IN2(n2592), .IN3(n2685), .Q(n2683) );
  INVX0 U2699 ( .INP(n2584), .ZN(n2685) );
  AO21X1 U2700 ( .IN1(n2686), .IN2(n2592), .IN3(n2684), .Q(n2584) );
  AO21X1 U2701 ( .IN1(N222), .IN2(N290), .IN3(n2687), .Q(n2686) );
  INVX0 U2702 ( .INP(n2688), .ZN(n2687) );
  NAND3X0 U2703 ( .IN1(N239), .IN2(n2688), .IN3(N273), .QN(n2592) );
  NAND3X0 U2704 ( .IN1(N239), .IN2(n2689), .IN3(N273), .QN(n2688) );
  NAND2X0 U2705 ( .IN1(N222), .IN2(N290), .QN(n2689) );
  XNOR2X1 U2706 ( .IN1(n2690), .IN2(keyinput33), .Q(n2680) );
  NAND2X0 U2707 ( .IN1(n2691), .IN2(n2692), .QN(n2690) );
  NAND2X0 U2708 ( .IN1(N103), .IN2(N409), .QN(n2635) );
  NAND2X0 U2709 ( .IN1(n2603), .IN2(n2693), .QN(N5672) );
  NAND3X0 U2710 ( .IN1(N494), .IN2(n2694), .IN3(N1), .QN(n2693) );
  AO21X1 U2711 ( .IN1(N1), .IN2(N494), .IN3(n2694), .Q(n2603) );
  NAND2X0 U2712 ( .IN1(n2604), .IN2(n2695), .QN(n2694) );
  NAND3X0 U2713 ( .IN1(n2696), .IN2(n2697), .IN3(n2698), .QN(n2695) );
  AO21X1 U2714 ( .IN1(n2696), .IN2(n2697), .IN3(n2698), .Q(n2604) );
  NAND2X0 U2715 ( .IN1(n2609), .IN2(n2699), .QN(n2698) );
  NAND3X0 U2716 ( .IN1(N477), .IN2(n2700), .IN3(N18), .QN(n2699) );
  AO21X1 U2717 ( .IN1(N18), .IN2(N477), .IN3(n2700), .Q(n2609) );
  NAND2X0 U2718 ( .IN1(n2610), .IN2(n2701), .QN(n2700) );
  NAND3X0 U2719 ( .IN1(n2702), .IN2(n2703), .IN3(n2704), .QN(n2701) );
  AO21X1 U2720 ( .IN1(n2704), .IN2(n2703), .IN3(n2702), .Q(n2610) );
  NAND2X0 U2721 ( .IN1(n2613), .IN2(n2705), .QN(n2702) );
  NAND3X0 U2722 ( .IN1(N460), .IN2(n2706), .IN3(N35), .QN(n2705) );
  AO21X1 U2723 ( .IN1(N35), .IN2(N460), .IN3(n2706), .Q(n2613) );
  NAND2X0 U2724 ( .IN1(n2614), .IN2(n2707), .QN(n2706) );
  NAND3X0 U2725 ( .IN1(n2708), .IN2(n2709), .IN3(n2710), .QN(n2707) );
  AO21X1 U2726 ( .IN1(n2708), .IN2(n2709), .IN3(n2710), .Q(n2614) );
  NAND2X0 U2727 ( .IN1(n2620), .IN2(n2711), .QN(n2710) );
  NAND3X0 U2728 ( .IN1(N443), .IN2(n2712), .IN3(N52), .QN(n2711) );
  AO21X1 U2729 ( .IN1(N52), .IN2(N443), .IN3(n2712), .Q(n2620) );
  NAND2X0 U2730 ( .IN1(n2621), .IN2(n2713), .QN(n2712) );
  NAND3X0 U2731 ( .IN1(n2714), .IN2(n2715), .IN3(n2716), .QN(n2713) );
  AO21X1 U2732 ( .IN1(n2714), .IN2(n2715), .IN3(n2716), .Q(n2621) );
  NAND2X0 U2733 ( .IN1(n2626), .IN2(n2717), .QN(n2716) );
  NAND3X0 U2734 ( .IN1(N426), .IN2(n2718), .IN3(N69), .QN(n2717) );
  AO21X1 U2735 ( .IN1(N69), .IN2(N426), .IN3(n2718), .Q(n2626) );
  NAND2X0 U2736 ( .IN1(n2627), .IN2(n2719), .QN(n2718) );
  NAND3X0 U2737 ( .IN1(n2720), .IN2(n2721), .IN3(n2722), .QN(n2719) );
  AO21X1 U2738 ( .IN1(n2722), .IN2(n2721), .IN3(n2720), .Q(n2627) );
  NAND2X0 U2739 ( .IN1(n2632), .IN2(n2723), .QN(n2720) );
  NAND3X0 U2740 ( .IN1(N409), .IN2(n2724), .IN3(N86), .QN(n2723) );
  AO21X1 U2741 ( .IN1(N86), .IN2(N409), .IN3(n2724), .Q(n2632) );
  XNOR2X1 U2742 ( .IN1(n2725), .IN2(keyinput70), .Q(n2724) );
  NAND2X0 U2743 ( .IN1(n2633), .IN2(n2726), .QN(n2725) );
  NAND3X0 U2744 ( .IN1(n2727), .IN2(n2728), .IN3(n2729), .QN(n2726) );
  AO21X1 U2745 ( .IN1(n2727), .IN2(n2728), .IN3(n2729), .Q(n2633) );
  NAND2X0 U2746 ( .IN1(n2642), .IN2(n2730), .QN(n2729) );
  NAND3X0 U2747 ( .IN1(N392), .IN2(n2731), .IN3(N103), .QN(n2730) );
  AO21X1 U2748 ( .IN1(N103), .IN2(N392), .IN3(n2731), .Q(n2642) );
  NAND2X0 U2749 ( .IN1(n2641), .IN2(n2732), .QN(n2731) );
  NAND4X0 U2750 ( .IN1(n2733), .IN2(n2734), .IN3(n2735), .IN4(n2736), .QN(
        n2732) );
  AO22X1 U2751 ( .IN1(n2735), .IN2(n2736), .IN3(n2733), .IN4(n2734), .Q(n2641)
         );
  AO21X1 U2752 ( .IN1(N120), .IN2(N375), .IN3(n2737), .Q(n2734) );
  INVX0 U2753 ( .INP(n2653), .ZN(n2737) );
  XOR2X1 U2754 ( .IN1(n2738), .IN2(keyinput54), .Q(n2733) );
  NAND2X0 U2755 ( .IN1(n2739), .IN2(n2653), .QN(n2738) );
  AO21X1 U2756 ( .IN1(N120), .IN2(N375), .IN3(n2740), .Q(n2653) );
  XOR2X1 U2757 ( .IN1(n2741), .IN2(keyinput50), .Q(n2740) );
  XNOR2X1 U2758 ( .IN1(keyinput50), .IN2(n2741), .Q(n2739) );
  XOR2X1 U2759 ( .IN1(n2651), .IN2(n2652), .Q(n2741) );
  NOR2X0 U2760 ( .IN1(n2742), .IN2(n2743), .QN(n2652) );
  INVX0 U2761 ( .INP(n2744), .ZN(n2743) );
  NAND2X0 U2762 ( .IN1(n2662), .IN2(n2745), .QN(n2651) );
  NAND3X0 U2763 ( .IN1(N358), .IN2(n2746), .IN3(N137), .QN(n2745) );
  AO21X1 U2764 ( .IN1(N137), .IN2(N358), .IN3(n2746), .Q(n2662) );
  NAND2X0 U2765 ( .IN1(n2663), .IN2(n2747), .QN(n2746) );
  NAND3X0 U2766 ( .IN1(n2748), .IN2(n2749), .IN3(n2750), .QN(n2747) );
  AO21X1 U2767 ( .IN1(n2748), .IN2(n2749), .IN3(n2750), .Q(n2663) );
  NAND2X0 U2768 ( .IN1(n2669), .IN2(n2751), .QN(n2750) );
  NAND3X0 U2769 ( .IN1(N154), .IN2(N341), .IN3(n2752), .QN(n2751) );
  AO21X1 U2770 ( .IN1(N154), .IN2(N341), .IN3(n2752), .Q(n2669) );
  XOR2X1 U2771 ( .IN1(n2753), .IN2(keyinput41), .Q(n2752) );
  NAND2X0 U2772 ( .IN1(n2670), .IN2(n2754), .QN(n2753) );
  NAND3X0 U2773 ( .IN1(n2755), .IN2(n2756), .IN3(n2757), .QN(n2754) );
  AO21X1 U2774 ( .IN1(n2755), .IN2(n2756), .IN3(n2757), .Q(n2670) );
  NAND2X0 U2775 ( .IN1(n2675), .IN2(n2758), .QN(n2757) );
  NAND3X0 U2776 ( .IN1(N324), .IN2(n2759), .IN3(N171), .QN(n2758) );
  AO21X1 U2777 ( .IN1(N171), .IN2(N324), .IN3(n2759), .Q(n2675) );
  NAND2X0 U2778 ( .IN1(n2676), .IN2(n2760), .QN(n2759) );
  NAND3X0 U2779 ( .IN1(n2761), .IN2(n2762), .IN3(n2763), .QN(n2760) );
  AO21X1 U2780 ( .IN1(n2761), .IN2(n2762), .IN3(n2763), .Q(n2676) );
  OAI21X1 U2781 ( .IN1(n2764), .IN2(n2765), .IN3(n2691), .QN(n2763) );
  XOR2X1 U2782 ( .IN1(n2766), .IN2(keyinput30), .Q(n2691) );
  NAND2X0 U2783 ( .IN1(n2764), .IN2(n2765), .QN(n2766) );
  NAND2X0 U2784 ( .IN1(N188), .IN2(N307), .QN(n2765) );
  AO21X1 U2785 ( .IN1(n2684), .IN2(n2692), .IN3(n2767), .Q(n2764) );
  XOR2X1 U2786 ( .IN1(keyinput29), .IN2(n2768), .Q(n2767) );
  NOR2X0 U2787 ( .IN1(n2769), .IN2(n2770), .QN(n2768) );
  INVX0 U2788 ( .INP(n2769), .ZN(n2692) );
  NOR2X0 U2789 ( .IN1(n2771), .IN2(n2770), .QN(n2769) );
  NOR3X0 U2790 ( .IN1(n2772), .IN2(n2773), .IN3(n2774), .QN(n2770) );
  AOI21X1 U2791 ( .IN1(n2775), .IN2(n2776), .IN3(n2684), .QN(n2771) );
  AND3X1 U2792 ( .IN1(N273), .IN2(n2775), .IN3(N222), .Q(n2684) );
  NAND3X0 U2793 ( .IN1(N273), .IN2(n2776), .IN3(N222), .QN(n2775) );
  NAND2X0 U2794 ( .IN1(N205), .IN2(N290), .QN(n2776) );
  INVX0 U2795 ( .INP(n2777), .ZN(n2704) );
  NOR2X0 U2796 ( .IN1(n2772), .IN2(n2601), .QN(N545) );
  NAND2X0 U2797 ( .IN1(n2696), .IN2(n2778), .QN(N5308) );
  NAND3X0 U2798 ( .IN1(N477), .IN2(n2779), .IN3(N1), .QN(n2778) );
  AO21X1 U2799 ( .IN1(N1), .IN2(N477), .IN3(n2779), .Q(n2696) );
  NAND2X0 U2800 ( .IN1(n2697), .IN2(n2780), .QN(n2779) );
  NAND3X0 U2801 ( .IN1(n2781), .IN2(n2782), .IN3(n2783), .QN(n2780) );
  AO21X1 U2802 ( .IN1(n2781), .IN2(n2782), .IN3(n2783), .Q(n2697) );
  NAND2X0 U2803 ( .IN1(n2703), .IN2(n2784), .QN(n2783) );
  NAND3X0 U2804 ( .IN1(N460), .IN2(n2785), .IN3(N18), .QN(n2784) );
  AO21X1 U2805 ( .IN1(N18), .IN2(N460), .IN3(n2785), .Q(n2703) );
  AO21X1 U2806 ( .IN1(n2786), .IN2(n2787), .IN3(n2777), .Q(n2785) );
  XOR2X1 U2807 ( .IN1(n2788), .IN2(keyinput95), .Q(n2777) );
  OR2X1 U2808 ( .IN1(n2787), .IN2(n2786), .Q(n2788) );
  NAND2X0 U2809 ( .IN1(n2708), .IN2(n2789), .QN(n2787) );
  NAND3X0 U2810 ( .IN1(N443), .IN2(n2790), .IN3(N35), .QN(n2789) );
  AO21X1 U2811 ( .IN1(N35), .IN2(N443), .IN3(n2790), .Q(n2708) );
  NAND2X0 U2812 ( .IN1(n2709), .IN2(n2791), .QN(n2790) );
  NAND3X0 U2813 ( .IN1(n2792), .IN2(n2793), .IN3(n2794), .QN(n2791) );
  AO21X1 U2814 ( .IN1(n2792), .IN2(n2793), .IN3(n2794), .Q(n2709) );
  NAND2X0 U2815 ( .IN1(n2714), .IN2(n2795), .QN(n2794) );
  NAND3X0 U2816 ( .IN1(N426), .IN2(n2796), .IN3(N52), .QN(n2795) );
  AO21X1 U2817 ( .IN1(N52), .IN2(N426), .IN3(n2796), .Q(n2714) );
  NAND2X0 U2818 ( .IN1(n2715), .IN2(n2797), .QN(n2796) );
  NAND3X0 U2819 ( .IN1(n2798), .IN2(n2799), .IN3(n2800), .QN(n2797) );
  AO21X1 U2820 ( .IN1(n2798), .IN2(n2799), .IN3(n2800), .Q(n2715) );
  NAND2X0 U2821 ( .IN1(n2721), .IN2(n2801), .QN(n2800) );
  NAND3X0 U2822 ( .IN1(N409), .IN2(n2802), .IN3(N69), .QN(n2801) );
  AO21X1 U2823 ( .IN1(N69), .IN2(N409), .IN3(n2802), .Q(n2721) );
  NAND2X0 U2824 ( .IN1(n2722), .IN2(n2803), .QN(n2802) );
  NAND3X0 U2825 ( .IN1(n2804), .IN2(n2805), .IN3(n2806), .QN(n2803) );
  XNOR2X1 U2826 ( .IN1(keyinput65), .IN2(n2807), .Q(n2722) );
  AOI21X1 U2827 ( .IN1(n2805), .IN2(n2804), .IN3(n2806), .QN(n2807) );
  OA22X1 U2828 ( .IN1(n2808), .IN2(n2809), .IN3(keyinput63), .IN4(n2810), .Q(
        n2806) );
  OA21X1 U2829 ( .IN1(n1975), .IN2(n2811), .IN3(n2727), .Q(n2810) );
  INVX0 U2830 ( .INP(n2808), .ZN(n2727) );
  NOR3X0 U2831 ( .IN1(n2812), .IN2(n2813), .IN3(n2814), .QN(n2809) );
  OA21X1 U2832 ( .IN1(n1975), .IN2(n2811), .IN3(keyinput63), .Q(n2814) );
  OA22X1 U2833 ( .IN1(n2811), .IN2(n1975), .IN3(n2812), .IN4(n2813), .Q(n2808)
         );
  AND2X1 U2834 ( .IN1(n2815), .IN2(n2728), .Q(n2813) );
  XOR2X1 U2835 ( .IN1(n2816), .IN2(keyinput59), .Q(n2812) );
  NAND2X0 U2836 ( .IN1(n2728), .IN2(n2817), .QN(n2816) );
  NAND2X0 U2837 ( .IN1(n2815), .IN2(n2817), .QN(n2728) );
  AND2X1 U2838 ( .IN1(n2735), .IN2(n2818), .Q(n2815) );
  NAND3X0 U2839 ( .IN1(N375), .IN2(n2819), .IN3(N103), .QN(n2818) );
  AO21X1 U2840 ( .IN1(N103), .IN2(N375), .IN3(n2819), .Q(n2735) );
  NAND2X0 U2841 ( .IN1(n2736), .IN2(n2820), .QN(n2819) );
  NAND3X0 U2842 ( .IN1(n2821), .IN2(n2822), .IN3(n2823), .QN(n2820) );
  AO21X1 U2843 ( .IN1(n2821), .IN2(n2822), .IN3(n2823), .Q(n2736) );
  AO21X1 U2844 ( .IN1(n2824), .IN2(n2825), .IN3(n2742), .Q(n2823) );
  XOR2X1 U2845 ( .IN1(n2826), .IN2(keyinput46), .Q(n2742) );
  OR2X1 U2846 ( .IN1(n2825), .IN2(n2824), .Q(n2826) );
  NAND2X0 U2847 ( .IN1(n2744), .IN2(n2827), .QN(n2825) );
  NAND3X0 U2848 ( .IN1(n2828), .IN2(n2829), .IN3(n2830), .QN(n2827) );
  AO21X1 U2849 ( .IN1(n2828), .IN2(n2829), .IN3(n2830), .Q(n2744) );
  NAND2X0 U2850 ( .IN1(n2748), .IN2(n2831), .QN(n2830) );
  NAND3X0 U2851 ( .IN1(N341), .IN2(n2832), .IN3(N137), .QN(n2831) );
  AO21X1 U2852 ( .IN1(N137), .IN2(N341), .IN3(n2832), .Q(n2748) );
  NAND2X0 U2853 ( .IN1(n2749), .IN2(n2833), .QN(n2832) );
  NAND3X0 U2854 ( .IN1(n2834), .IN2(n2835), .IN3(n2836), .QN(n2833) );
  AO21X1 U2855 ( .IN1(n2834), .IN2(n2835), .IN3(n2836), .Q(n2749) );
  XNOR2X1 U2856 ( .IN1(n2837), .IN2(keyinput38), .Q(n2836) );
  NAND2X0 U2857 ( .IN1(n2755), .IN2(n2838), .QN(n2837) );
  NAND3X0 U2858 ( .IN1(N324), .IN2(n2839), .IN3(N154), .QN(n2838) );
  AO21X1 U2859 ( .IN1(N154), .IN2(N324), .IN3(n2839), .Q(n2755) );
  NAND2X0 U2860 ( .IN1(n2756), .IN2(n2840), .QN(n2839) );
  NAND3X0 U2861 ( .IN1(n2841), .IN2(n2842), .IN3(n2843), .QN(n2840) );
  AO21X1 U2862 ( .IN1(n2843), .IN2(n2842), .IN3(n2841), .Q(n2756) );
  NAND2X0 U2863 ( .IN1(n2761), .IN2(n2844), .QN(n2841) );
  NAND4X0 U2864 ( .IN1(n2845), .IN2(N171), .IN3(N307), .IN4(n2846), .QN(n2844)
         );
  AO22X1 U2865 ( .IN1(N171), .IN2(N307), .IN3(n2845), .IN4(n2846), .Q(n2761)
         );
  NAND2X0 U2866 ( .IN1(n2847), .IN2(n2762), .QN(n2846) );
  XOR2X1 U2867 ( .IN1(n2848), .IN2(keyinput28), .Q(n2845) );
  NAND2X0 U2868 ( .IN1(n2849), .IN2(n2762), .QN(n2848) );
  NAND2X0 U2869 ( .IN1(n2849), .IN2(n2847), .QN(n2762) );
  AOI21X1 U2870 ( .IN1(n2850), .IN2(n2851), .IN3(n2773), .QN(n2849) );
  NOR2X0 U2871 ( .IN1(n2851), .IN2(n2850), .QN(n2773) );
  AND2X1 U2872 ( .IN1(N188), .IN2(N290), .Q(n2851) );
  OA21X1 U2873 ( .IN1(n2772), .IN2(n2774), .IN3(keyinput23), .Q(n2850) );
  INVX0 U2874 ( .INP(N205), .ZN(n2774) );
  INVX0 U2875 ( .INP(N273), .ZN(n2772) );
  NOR2X0 U2876 ( .IN1(n2000), .IN2(n2131), .QN(n2824) );
  INVX0 U2877 ( .INP(N358), .ZN(n2131) );
  INVX0 U2878 ( .INP(N392), .ZN(n1975) );
  INVX0 U2879 ( .INP(N86), .ZN(n2811) );
  AND2X1 U2880 ( .IN1(n2852), .IN2(n2853), .Q(n2786) );
  AO21X1 U2881 ( .IN1(n2854), .IN2(n2855), .IN3(n2856), .Q(n2852) );
  NAND2X0 U2882 ( .IN1(n2781), .IN2(n2857), .QN(N4946) );
  NAND3X0 U2883 ( .IN1(N1), .IN2(N460), .IN3(n2858), .QN(n2857) );
  AO21X1 U2884 ( .IN1(N1), .IN2(N460), .IN3(n2858), .Q(n2781) );
  AND2X1 U2885 ( .IN1(n2859), .IN2(n2860), .Q(n2858) );
  AO21X1 U2886 ( .IN1(n2861), .IN2(n2862), .IN3(n2863), .Q(n2860) );
  INVX0 U2887 ( .INP(n2782), .ZN(n2863) );
  XOR2X1 U2888 ( .IN1(n2864), .IN2(keyinput97), .Q(n2859) );
  NAND3X0 U2889 ( .IN1(n2865), .IN2(n2853), .IN3(n2782), .QN(n2864) );
  NAND3X0 U2890 ( .IN1(n2865), .IN2(n2853), .IN3(n2866), .QN(n2782) );
  NAND2X0 U2891 ( .IN1(n2861), .IN2(n2862), .QN(n2866) );
  AO21X1 U2892 ( .IN1(N18), .IN2(N443), .IN3(n2867), .Q(n2853) );
  NAND3X0 U2893 ( .IN1(N443), .IN2(n2867), .IN3(N18), .QN(n2865) );
  XNOR2X1 U2894 ( .IN1(n2856), .IN2(n2868), .Q(n2867) );
  AND2X1 U2895 ( .IN1(n2854), .IN2(n2855), .Q(n2868) );
  NAND2X0 U2896 ( .IN1(n2869), .IN2(n2870), .QN(n2854) );
  INVX0 U2897 ( .INP(n2871), .ZN(n2869) );
  NAND2X0 U2898 ( .IN1(n2792), .IN2(n2872), .QN(n2856) );
  NAND3X0 U2899 ( .IN1(N426), .IN2(n2873), .IN3(N35), .QN(n2872) );
  AO21X1 U2900 ( .IN1(N35), .IN2(N426), .IN3(n2873), .Q(n2792) );
  NAND2X0 U2901 ( .IN1(n2793), .IN2(n2874), .QN(n2873) );
  NAND3X0 U2902 ( .IN1(n2875), .IN2(n2876), .IN3(n2877), .QN(n2874) );
  AO21X1 U2903 ( .IN1(n2877), .IN2(n2876), .IN3(n2875), .Q(n2793) );
  NAND2X0 U2904 ( .IN1(n2798), .IN2(n2878), .QN(n2875) );
  NAND4X0 U2905 ( .IN1(N52), .IN2(N409), .IN3(n2879), .IN4(n2880), .QN(n2878)
         );
  AO22X1 U2906 ( .IN1(N52), .IN2(N409), .IN3(n2879), .IN4(n2880), .Q(n2798) );
  NAND2X0 U2907 ( .IN1(n2881), .IN2(n2799), .QN(n2880) );
  XNOR2X1 U2908 ( .IN1(n2882), .IN2(keyinput68), .Q(n2879) );
  NAND2X0 U2909 ( .IN1(n2883), .IN2(n2799), .QN(n2882) );
  NAND2X0 U2910 ( .IN1(n2881), .IN2(n2883), .QN(n2799) );
  AND2X1 U2911 ( .IN1(n2804), .IN2(n2884), .Q(n2881) );
  NAND3X0 U2912 ( .IN1(N392), .IN2(n2885), .IN3(N69), .QN(n2884) );
  AO21X1 U2913 ( .IN1(N69), .IN2(N392), .IN3(n2885), .Q(n2804) );
  NAND2X0 U2914 ( .IN1(n2805), .IN2(n2886), .QN(n2885) );
  NAND4X0 U2915 ( .IN1(n2887), .IN2(n2888), .IN3(n2889), .IN4(n2890), .QN(
        n2886) );
  AO22X1 U2916 ( .IN1(n2887), .IN2(n2888), .IN3(n2889), .IN4(n2890), .Q(n2805)
         );
  NAND2X0 U2917 ( .IN1(n2891), .IN2(n2892), .QN(n2888) );
  INVX0 U2918 ( .INP(n2817), .ZN(n2891) );
  NAND2X0 U2919 ( .IN1(n2893), .IN2(n2894), .QN(n2817) );
  XOR2X1 U2920 ( .IN1(n2895), .IN2(keyinput53), .Q(n2887) );
  NAND2X0 U2921 ( .IN1(n2894), .IN2(n2896), .QN(n2895) );
  NAND3X0 U2922 ( .IN1(n2896), .IN2(n2892), .IN3(n2893), .QN(n2894) );
  XNOR2X1 U2923 ( .IN1(keyinput49), .IN2(n2897), .Q(n2893) );
  AOI21X1 U2924 ( .IN1(n2898), .IN2(n2899), .IN3(n2900), .QN(n2897) );
  NAND3X0 U2925 ( .IN1(n2899), .IN2(n2898), .IN3(n2900), .QN(n2892) );
  NAND2X0 U2926 ( .IN1(n2821), .IN2(n2901), .QN(n2900) );
  NAND3X0 U2927 ( .IN1(N358), .IN2(n2902), .IN3(N103), .QN(n2901) );
  AO21X1 U2928 ( .IN1(N103), .IN2(N358), .IN3(n2902), .Q(n2821) );
  NAND2X0 U2929 ( .IN1(n2822), .IN2(n2903), .QN(n2902) );
  NAND3X0 U2930 ( .IN1(n2904), .IN2(n2905), .IN3(n2906), .QN(n2903) );
  AO21X1 U2931 ( .IN1(n2904), .IN2(n2905), .IN3(n2906), .Q(n2822) );
  NAND2X0 U2932 ( .IN1(n2828), .IN2(n2907), .QN(n2906) );
  NAND3X0 U2933 ( .IN1(N341), .IN2(n2908), .IN3(N120), .QN(n2907) );
  AO21X1 U2934 ( .IN1(N120), .IN2(N341), .IN3(n2908), .Q(n2828) );
  NAND2X0 U2935 ( .IN1(n2829), .IN2(n2909), .QN(n2908) );
  NAND3X0 U2936 ( .IN1(n2910), .IN2(n2911), .IN3(n2912), .QN(n2909) );
  AO21X1 U2937 ( .IN1(n2910), .IN2(n2911), .IN3(n2912), .Q(n2829) );
  NAND2X0 U2938 ( .IN1(n2834), .IN2(n2913), .QN(n2912) );
  NAND3X0 U2939 ( .IN1(N324), .IN2(n2914), .IN3(N137), .QN(n2913) );
  AO21X1 U2940 ( .IN1(N137), .IN2(N324), .IN3(n2914), .Q(n2834) );
  NAND2X0 U2941 ( .IN1(n2835), .IN2(n2915), .QN(n2914) );
  NAND3X0 U2942 ( .IN1(n2916), .IN2(n2917), .IN3(n2918), .QN(n2915) );
  AO21X1 U2943 ( .IN1(n2916), .IN2(n2917), .IN3(n2918), .Q(n2835) );
  NAND2X0 U2944 ( .IN1(n2842), .IN2(n2919), .QN(n2918) );
  NAND3X0 U2945 ( .IN1(N307), .IN2(n2920), .IN3(N154), .QN(n2919) );
  AO21X1 U2946 ( .IN1(N154), .IN2(N307), .IN3(n2920), .Q(n2842) );
  OAI21X1 U2947 ( .IN1(n2921), .IN2(n2922), .IN3(n2843), .QN(n2920) );
  XNOR2X1 U2948 ( .IN1(keyinput26), .IN2(n2923), .Q(n2843) );
  OA21X1 U2949 ( .IN1(n2924), .IN2(n2922), .IN3(n2921), .Q(n2923) );
  OA21X1 U2950 ( .IN1(n2925), .IN2(n2926), .IN3(n2927), .Q(n2924) );
  INVX0 U2951 ( .INP(N171), .ZN(n2926) );
  INVX0 U2952 ( .INP(n2847), .ZN(n2922) );
  NAND3X0 U2953 ( .IN1(N273), .IN2(n2927), .IN3(N188), .QN(n2847) );
  NAND3X0 U2954 ( .IN1(N273), .IN2(n2928), .IN3(N188), .QN(n2927) );
  NAND2X0 U2955 ( .IN1(N171), .IN2(N290), .QN(n2928) );
  NAND2X0 U2956 ( .IN1(N86), .IN2(N375), .QN(n2896) );
  AO22X1 U2957 ( .IN1(n2929), .IN2(n2930), .IN3(n2931), .IN4(n2932), .Q(n2883)
         );
  NAND2X0 U2958 ( .IN1(n2861), .IN2(n2933), .QN(N4591) );
  NAND3X0 U2959 ( .IN1(N443), .IN2(n2934), .IN3(N1), .QN(n2933) );
  AO21X1 U2960 ( .IN1(N1), .IN2(N443), .IN3(n2934), .Q(n2861) );
  NAND2X0 U2961 ( .IN1(n2862), .IN2(n2935), .QN(n2934) );
  NAND3X0 U2962 ( .IN1(n2936), .IN2(n2937), .IN3(n2938), .QN(n2935) );
  AO21X1 U2963 ( .IN1(n2936), .IN2(n2937), .IN3(n2938), .Q(n2862) );
  NAND2X0 U2964 ( .IN1(n2855), .IN2(n2939), .QN(n2938) );
  NAND4X0 U2965 ( .IN1(N18), .IN2(N426), .IN3(n2940), .IN4(n2941), .QN(n2939)
         );
  AO22X1 U2966 ( .IN1(N18), .IN2(N426), .IN3(n2940), .IN4(n2941), .Q(n2855) );
  OR2X1 U2967 ( .IN1(n2870), .IN2(n2871), .Q(n2941) );
  XNOR2X1 U2968 ( .IN1(n2942), .IN2(keyinput78), .Q(n2940) );
  NAND2X0 U2969 ( .IN1(n2871), .IN2(n2870), .QN(n2942) );
  AO22X1 U2970 ( .IN1(n2943), .IN2(n2944), .IN3(n2945), .IN4(n2946), .Q(n2870)
         );
  XOR2X1 U2971 ( .IN1(keyinput75), .IN2(n2947), .Q(n2871) );
  OA21X1 U2972 ( .IN1(n2948), .IN2(n2949), .IN3(n2877), .Q(n2947) );
  XNOR2X1 U2973 ( .IN1(n2950), .IN2(keyinput71), .Q(n2877) );
  NAND2X0 U2974 ( .IN1(n2948), .IN2(n2949), .QN(n2950) );
  NAND2X0 U2975 ( .IN1(N35), .IN2(N409), .QN(n2949) );
  AND2X1 U2976 ( .IN1(n2951), .IN2(n2876), .Q(n2948) );
  AO21X1 U2977 ( .IN1(n2952), .IN2(n2953), .IN3(n2954), .Q(n2876) );
  NAND3X0 U2978 ( .IN1(n2952), .IN2(n2953), .IN3(n2954), .QN(n2951) );
  XNOR2X1 U2979 ( .IN1(n2930), .IN2(n2929), .Q(n2954) );
  XOR2X1 U2980 ( .IN1(n2931), .IN2(n2932), .Q(n2929) );
  NAND2X0 U2981 ( .IN1(n2955), .IN2(n2956), .QN(n2932) );
  INVX0 U2982 ( .INP(n2957), .ZN(n2956) );
  AND2X1 U2983 ( .IN1(n2889), .IN2(n2958), .Q(n2931) );
  NAND3X0 U2984 ( .IN1(N375), .IN2(n2959), .IN3(N69), .QN(n2958) );
  AO21X1 U2985 ( .IN1(N69), .IN2(N375), .IN3(n2959), .Q(n2889) );
  NAND2X0 U2986 ( .IN1(n2890), .IN2(n2960), .QN(n2959) );
  NAND3X0 U2987 ( .IN1(n2961), .IN2(n2962), .IN3(n2963), .QN(n2960) );
  AO21X1 U2988 ( .IN1(n2961), .IN2(n2962), .IN3(n2963), .Q(n2890) );
  NAND2X0 U2989 ( .IN1(n2899), .IN2(n2964), .QN(n2963) );
  NAND3X0 U2990 ( .IN1(N358), .IN2(n2965), .IN3(N86), .QN(n2964) );
  AO21X1 U2991 ( .IN1(N86), .IN2(N358), .IN3(n2965), .Q(n2899) );
  NAND2X0 U2992 ( .IN1(n2898), .IN2(n2966), .QN(n2965) );
  NAND3X0 U2993 ( .IN1(n2967), .IN2(n2968), .IN3(n2969), .QN(n2966) );
  AO21X1 U2994 ( .IN1(n2967), .IN2(n2968), .IN3(n2969), .Q(n2898) );
  NAND2X0 U2995 ( .IN1(n2904), .IN2(n2970), .QN(n2969) );
  NAND3X0 U2996 ( .IN1(N341), .IN2(n2971), .IN3(N103), .QN(n2970) );
  AO21X1 U2997 ( .IN1(N103), .IN2(N341), .IN3(n2971), .Q(n2904) );
  NAND2X0 U2998 ( .IN1(n2905), .IN2(n2972), .QN(n2971) );
  NAND3X0 U2999 ( .IN1(n2973), .IN2(n2974), .IN3(n2975), .QN(n2972) );
  AO21X1 U3000 ( .IN1(n2973), .IN2(n2974), .IN3(n2975), .Q(n2905) );
  NAND2X0 U3001 ( .IN1(n2910), .IN2(n2976), .QN(n2975) );
  NAND3X0 U3002 ( .IN1(N324), .IN2(n2977), .IN3(N120), .QN(n2976) );
  AO21X1 U3003 ( .IN1(N120), .IN2(N324), .IN3(n2977), .Q(n2910) );
  NAND2X0 U3004 ( .IN1(n2911), .IN2(n2978), .QN(n2977) );
  NAND3X0 U3005 ( .IN1(n2979), .IN2(n2980), .IN3(n2981), .QN(n2978) );
  AO21X1 U3006 ( .IN1(n2979), .IN2(n2980), .IN3(n2981), .Q(n2911) );
  NAND2X0 U3007 ( .IN1(n2916), .IN2(n2982), .QN(n2981) );
  NAND3X0 U3008 ( .IN1(N307), .IN2(n2983), .IN3(N137), .QN(n2982) );
  AO21X1 U3009 ( .IN1(N137), .IN2(N307), .IN3(n2983), .Q(n2916) );
  AO21X1 U3010 ( .IN1(n2984), .IN2(n2921), .IN3(n2985), .Q(n2983) );
  INVX0 U3011 ( .INP(n2917), .ZN(n2985) );
  AO21X1 U3012 ( .IN1(n2986), .IN2(n2921), .IN3(n2984), .Q(n2917) );
  OAI21X1 U3013 ( .IN1(n1907), .IN2(n2925), .IN3(n2987), .QN(n2986) );
  INVX0 U3014 ( .INP(N154), .ZN(n1907) );
  NAND3X0 U3015 ( .IN1(N273), .IN2(n2987), .IN3(N171), .QN(n2921) );
  NAND3X0 U3016 ( .IN1(N273), .IN2(n2988), .IN3(N171), .QN(n2987) );
  NAND2X0 U3017 ( .IN1(N154), .IN2(N290), .QN(n2988) );
  INVX0 U3018 ( .INP(n2989), .ZN(n2984) );
  INVX0 U3019 ( .INP(n2990), .ZN(n2980) );
  XNOR2X1 U3020 ( .IN1(n2991), .IN2(keyinput6), .Q(n2930) );
  NAND2X0 U3021 ( .IN1(N52), .IN2(N392), .QN(n2991) );
  OA21X1 U3022 ( .IN1(n2992), .IN2(n2993), .IN3(n2994), .Q(N4241) );
  XOR2X1 U3023 ( .IN1(n2995), .IN2(keyinput85), .Q(n2994) );
  NAND2X0 U3024 ( .IN1(n2937), .IN2(n2996), .QN(n2995) );
  INVX0 U3025 ( .INP(n2937), .ZN(n2992) );
  NAND2X0 U3026 ( .IN1(n2997), .IN2(n2996), .QN(n2937) );
  NAND2X0 U3027 ( .IN1(N1), .IN2(N426), .QN(n2996) );
  INVX0 U3028 ( .INP(n2993), .ZN(n2997) );
  NAND2X0 U3029 ( .IN1(n2936), .IN2(n2998), .QN(n2993) );
  NAND3X0 U3030 ( .IN1(n2999), .IN2(n3000), .IN3(n3001), .QN(n2998) );
  AO21X1 U3031 ( .IN1(n2999), .IN2(n3000), .IN3(n3001), .Q(n2936) );
  XNOR2X1 U3032 ( .IN1(n2945), .IN2(n2946), .Q(n3001) );
  NAND2X0 U3033 ( .IN1(N18), .IN2(N409), .QN(n2946) );
  XOR2X1 U3034 ( .IN1(n2943), .IN2(n2944), .Q(n2945) );
  XOR2X1 U3035 ( .IN1(keyinput62), .IN2(n3002), .Q(n2944) );
  OA22X1 U3036 ( .IN1(n3003), .IN2(n3004), .IN3(n3005), .IN4(n3006), .Q(n3002)
         );
  OA21X1 U3037 ( .IN1(n3007), .IN2(n3008), .IN3(n2952), .Q(n2943) );
  XNOR2X1 U3038 ( .IN1(n3009), .IN2(keyinput61), .Q(n2952) );
  NAND2X0 U3039 ( .IN1(n3008), .IN2(n3007), .QN(n3009) );
  AND2X1 U3040 ( .IN1(n3010), .IN2(n2953), .Q(n3008) );
  AO221X1 U3041 ( .IN1(n3011), .IN2(n3012), .IN3(n3013), .IN4(n3014), .IN5(
        n2957), .Q(n2953) );
  NOR2X0 U3042 ( .IN1(n3012), .IN2(n3011), .QN(n2957) );
  NAND3X0 U3043 ( .IN1(n3013), .IN2(n3014), .IN3(n3015), .QN(n3010) );
  XNOR2X1 U3044 ( .IN1(n3012), .IN2(n3011), .Q(n3015) );
  XOR2X1 U3045 ( .IN1(n3016), .IN2(keyinput5), .Q(n3011) );
  NAND2X0 U3046 ( .IN1(N52), .IN2(N375), .QN(n3016) );
  NAND2X0 U3047 ( .IN1(n2955), .IN2(n3017), .QN(n3012) );
  NAND3X0 U3048 ( .IN1(n3018), .IN2(n3019), .IN3(n3020), .QN(n3017) );
  AO21X1 U3049 ( .IN1(n3018), .IN2(n3019), .IN3(n3020), .Q(n2955) );
  NAND2X0 U3050 ( .IN1(n2961), .IN2(n3021), .QN(n3020) );
  NAND3X0 U3051 ( .IN1(N358), .IN2(n3022), .IN3(N69), .QN(n3021) );
  AO21X1 U3052 ( .IN1(N69), .IN2(N358), .IN3(n3022), .Q(n2961) );
  NAND2X0 U3053 ( .IN1(n2962), .IN2(n3023), .QN(n3022) );
  NAND3X0 U3054 ( .IN1(n3024), .IN2(n3025), .IN3(n3026), .QN(n3023) );
  AO21X1 U3055 ( .IN1(n3026), .IN2(n3025), .IN3(n3024), .Q(n2962) );
  NAND2X0 U3056 ( .IN1(n2967), .IN2(n3027), .QN(n3024) );
  NAND3X0 U3057 ( .IN1(N341), .IN2(n3028), .IN3(N86), .QN(n3027) );
  AO21X1 U3058 ( .IN1(N86), .IN2(N341), .IN3(n3028), .Q(n2967) );
  NAND2X0 U3059 ( .IN1(n2968), .IN2(n3029), .QN(n3028) );
  NAND3X0 U3060 ( .IN1(n3030), .IN2(n3031), .IN3(n3032), .QN(n3029) );
  AO21X1 U3061 ( .IN1(n3030), .IN2(n3031), .IN3(n3032), .Q(n2968) );
  NAND2X0 U3062 ( .IN1(n2973), .IN2(n3033), .QN(n3032) );
  NAND3X0 U3063 ( .IN1(N324), .IN2(n3034), .IN3(N103), .QN(n3033) );
  AO21X1 U3064 ( .IN1(N103), .IN2(N324), .IN3(n3034), .Q(n2973) );
  NAND2X0 U3065 ( .IN1(n2974), .IN2(n3035), .QN(n3034) );
  NAND3X0 U3066 ( .IN1(n3036), .IN2(n3037), .IN3(n3038), .QN(n3035) );
  AO21X1 U3067 ( .IN1(n3036), .IN2(n3037), .IN3(n3038), .Q(n2974) );
  NAND2X0 U3068 ( .IN1(n2979), .IN2(n3039), .QN(n3038) );
  NAND3X0 U3069 ( .IN1(N307), .IN2(n3040), .IN3(N120), .QN(n3039) );
  AO21X1 U3070 ( .IN1(N120), .IN2(N307), .IN3(n3040), .Q(n2979) );
  AO21X1 U3071 ( .IN1(n3041), .IN2(n3042), .IN3(n2990), .Q(n3040) );
  NOR2X0 U3072 ( .IN1(n3042), .IN2(n3041), .QN(n2990) );
  XNOR2X1 U3073 ( .IN1(n3043), .IN2(keyinput25), .Q(n3042) );
  AND2X1 U3074 ( .IN1(n3044), .IN2(n2989), .Q(n3041) );
  NAND3X0 U3075 ( .IN1(N273), .IN2(n3045), .IN3(N154), .QN(n2989) );
  AO21X1 U3076 ( .IN1(N137), .IN2(N290), .IN3(n3046), .Q(n3044) );
  INVX0 U3077 ( .INP(n3045), .ZN(n3046) );
  NAND3X0 U3078 ( .IN1(N273), .IN2(n3047), .IN3(N154), .QN(n3045) );
  NAND2X0 U3079 ( .IN1(N137), .IN2(N290), .QN(n3047) );
  NAND2X0 U3080 ( .IN1(N35), .IN2(N392), .QN(n3007) );
  NAND2X0 U3081 ( .IN1(n2999), .IN2(n3048), .QN(N3895) );
  NAND3X0 U3082 ( .IN1(N409), .IN2(n3049), .IN3(N1), .QN(n3048) );
  AO21X1 U3083 ( .IN1(N1), .IN2(N409), .IN3(n3049), .Q(n2999) );
  NAND2X0 U3084 ( .IN1(n3000), .IN2(n3050), .QN(n3049) );
  NAND3X0 U3085 ( .IN1(n3051), .IN2(n3052), .IN3(n3053), .QN(n3050) );
  AO21X1 U3086 ( .IN1(n3051), .IN2(n3052), .IN3(n3053), .Q(n3000) );
  XNOR2X1 U3087 ( .IN1(n3005), .IN2(n3006), .Q(n3053) );
  XNOR2X1 U3088 ( .IN1(n3003), .IN2(n3004), .Q(n3006) );
  NAND2X0 U3089 ( .IN1(n3013), .IN2(n3054), .QN(n3004) );
  NAND3X0 U3090 ( .IN1(N375), .IN2(n3055), .IN3(N35), .QN(n3054) );
  AO21X1 U3091 ( .IN1(N35), .IN2(N375), .IN3(n3055), .Q(n3013) );
  NAND2X0 U3092 ( .IN1(n3014), .IN2(n3056), .QN(n3055) );
  NAND3X0 U3093 ( .IN1(n3057), .IN2(n3058), .IN3(n3059), .QN(n3056) );
  AO21X1 U3094 ( .IN1(n3057), .IN2(n3058), .IN3(n3059), .Q(n3014) );
  NAND2X0 U3095 ( .IN1(n3018), .IN2(n3060), .QN(n3059) );
  NAND3X0 U3096 ( .IN1(N358), .IN2(n3061), .IN3(N52), .QN(n3060) );
  AO21X1 U3097 ( .IN1(N52), .IN2(N358), .IN3(n3061), .Q(n3018) );
  NAND2X0 U3098 ( .IN1(n3019), .IN2(n3062), .QN(n3061) );
  NAND3X0 U3099 ( .IN1(n3063), .IN2(n3064), .IN3(n3065), .QN(n3062) );
  AO21X1 U3100 ( .IN1(n3065), .IN2(n3064), .IN3(n3063), .Q(n3019) );
  NAND2X0 U3101 ( .IN1(n3025), .IN2(n3066), .QN(n3063) );
  NAND3X0 U3102 ( .IN1(N341), .IN2(n3067), .IN3(N69), .QN(n3066) );
  AO21X1 U3103 ( .IN1(N69), .IN2(N341), .IN3(n3067), .Q(n3025) );
  NAND2X0 U3104 ( .IN1(n3026), .IN2(n3068), .QN(n3067) );
  NAND3X0 U3105 ( .IN1(n3069), .IN2(n3070), .IN3(n3071), .QN(n3068) );
  XOR2X1 U3106 ( .IN1(keyinput39), .IN2(n3072), .Q(n3026) );
  AOI21X1 U3107 ( .IN1(n3070), .IN2(n3071), .IN3(n3069), .QN(n3072) );
  NAND2X0 U3108 ( .IN1(n3030), .IN2(n3073), .QN(n3069) );
  NAND3X0 U3109 ( .IN1(N86), .IN2(N324), .IN3(n3074), .QN(n3073) );
  AO21X1 U3110 ( .IN1(N86), .IN2(N324), .IN3(n3074), .Q(n3030) );
  XOR2X1 U3111 ( .IN1(n3075), .IN2(keyinput35), .Q(n3074) );
  NAND2X0 U3112 ( .IN1(n3031), .IN2(n3076), .QN(n3075) );
  NAND3X0 U3113 ( .IN1(n3077), .IN2(n3078), .IN3(n3079), .QN(n3076) );
  AO21X1 U3114 ( .IN1(n3077), .IN2(n3078), .IN3(n3079), .Q(n3031) );
  NAND2X0 U3115 ( .IN1(n3036), .IN2(n3080), .QN(n3079) );
  NAND3X0 U3116 ( .IN1(N307), .IN2(n3081), .IN3(N103), .QN(n3080) );
  AO21X1 U3117 ( .IN1(N103), .IN2(N307), .IN3(n3081), .Q(n3036) );
  NAND2X0 U3118 ( .IN1(n3037), .IN2(n3082), .QN(n3081) );
  NAND4X0 U3119 ( .IN1(n3083), .IN2(n3084), .IN3(n3085), .IN4(n3043), .QN(
        n3082) );
  NAND2X0 U3120 ( .IN1(n2000), .IN2(n3086), .QN(n3085) );
  AO22X1 U3121 ( .IN1(n3084), .IN2(n3083), .IN3(n3087), .IN4(n3043), .Q(n3037)
         );
  NAND3X0 U3122 ( .IN1(N273), .IN2(n3086), .IN3(N137), .QN(n3043) );
  OAI21X1 U3123 ( .IN1(n2000), .IN2(n2925), .IN3(n3086), .QN(n3087) );
  NAND3X0 U3124 ( .IN1(N273), .IN2(n3088), .IN3(N137), .QN(n3086) );
  NAND2X0 U3125 ( .IN1(N120), .IN2(N290), .QN(n3088) );
  INVX0 U3126 ( .INP(N120), .ZN(n2000) );
  INVX0 U3127 ( .INP(n3089), .ZN(n3071) );
  INVX0 U3128 ( .INP(n3090), .ZN(n3070) );
  INVX0 U3129 ( .INP(n3091), .ZN(n3065) );
  AND2X1 U3130 ( .IN1(n3092), .IN2(n3093), .Q(n3003) );
  XOR2X1 U3131 ( .IN1(n3094), .IN2(keyinput3), .Q(n3005) );
  NAND2X0 U3132 ( .IN1(N18), .IN2(N392), .QN(n3094) );
  NAND2X0 U3133 ( .IN1(n3051), .IN2(n3095), .QN(N3552) );
  NAND3X0 U3134 ( .IN1(n3096), .IN2(n3097), .IN3(n3098), .QN(n3095) );
  AO21X1 U3135 ( .IN1(n3096), .IN2(n3097), .IN3(n3098), .Q(n3051) );
  XNOR2X1 U3136 ( .IN1(n3099), .IN2(keyinput1), .Q(n3098) );
  NAND2X0 U3137 ( .IN1(N1), .IN2(N392), .QN(n3099) );
  NAND2X0 U3138 ( .IN1(n3100), .IN2(n3052), .QN(n3097) );
  XOR2X1 U3139 ( .IN1(keyinput58), .IN2(n3101), .Q(n3096) );
  OA21X1 U3140 ( .IN1(n3102), .IN2(n3103), .IN3(n3052), .Q(n3101) );
  OAI21X1 U3141 ( .IN1(n3103), .IN2(n3102), .IN3(n3100), .QN(n3052) );
  AND2X1 U3142 ( .IN1(n3093), .IN2(n3104), .Q(n3100) );
  NAND3X0 U3143 ( .IN1(N375), .IN2(n3105), .IN3(N18), .QN(n3104) );
  AO21X1 U3144 ( .IN1(N18), .IN2(N375), .IN3(n3105), .Q(n3093) );
  NAND2X0 U3145 ( .IN1(n3092), .IN2(n3106), .QN(n3105) );
  NAND3X0 U3146 ( .IN1(n3107), .IN2(n3108), .IN3(n3109), .QN(n3106) );
  AO21X1 U3147 ( .IN1(n3107), .IN2(n3108), .IN3(n3109), .Q(n3092) );
  NAND2X0 U3148 ( .IN1(n3057), .IN2(n3110), .QN(n3109) );
  NAND3X0 U3149 ( .IN1(N35), .IN2(N358), .IN3(n3111), .QN(n3110) );
  AO21X1 U3150 ( .IN1(N35), .IN2(N358), .IN3(n3111), .Q(n3057) );
  XOR2X1 U3151 ( .IN1(n3112), .IN2(keyinput45), .Q(n3111) );
  NAND2X0 U3152 ( .IN1(n3058), .IN2(n3113), .QN(n3112) );
  NAND3X0 U3153 ( .IN1(n3114), .IN2(n3115), .IN3(n3116), .QN(n3113) );
  AO21X1 U3154 ( .IN1(n3114), .IN2(n3115), .IN3(n3116), .Q(n3058) );
  AO21X1 U3155 ( .IN1(n3117), .IN2(n3118), .IN3(n3091), .Q(n3116) );
  NOR2X0 U3156 ( .IN1(n3118), .IN2(n3117), .QN(n3091) );
  NAND2X0 U3157 ( .IN1(n3064), .IN2(n3119), .QN(n3118) );
  NAND3X0 U3158 ( .IN1(n3120), .IN2(n3121), .IN3(n3122), .QN(n3119) );
  AO21X1 U3159 ( .IN1(n3120), .IN2(n3121), .IN3(n3122), .Q(n3064) );
  AO21X1 U3160 ( .IN1(n3123), .IN2(n3124), .IN3(n3089), .Q(n3122) );
  XOR2X1 U3161 ( .IN1(n3125), .IN2(keyinput36), .Q(n3089) );
  OR2X1 U3162 ( .IN1(n3124), .IN2(n3123), .Q(n3125) );
  AO21X1 U3163 ( .IN1(n3126), .IN2(n3127), .IN3(n3090), .Q(n3124) );
  NOR2X0 U3164 ( .IN1(n3127), .IN2(n3126), .QN(n3090) );
  NAND2X0 U3165 ( .IN1(n3077), .IN2(n3128), .QN(n3127) );
  NAND3X0 U3166 ( .IN1(N307), .IN2(n3129), .IN3(N86), .QN(n3128) );
  AO21X1 U3167 ( .IN1(N86), .IN2(N307), .IN3(n3129), .Q(n3077) );
  NAND2X0 U3168 ( .IN1(n3078), .IN2(n3130), .QN(n3129) );
  NAND3X0 U3169 ( .IN1(n3131), .IN2(n3132), .IN3(n3133), .QN(n3130) );
  AO21X1 U3170 ( .IN1(n3131), .IN2(n3132), .IN3(n3133), .Q(n3078) );
  XOR2X1 U3171 ( .IN1(n3083), .IN2(n3084), .Q(n3133) );
  AND2X1 U3172 ( .IN1(N103), .IN2(N290), .Q(n3084) );
  XOR2X1 U3173 ( .IN1(n3134), .IN2(keyinput10), .Q(n3083) );
  NAND2X0 U3174 ( .IN1(N120), .IN2(N273), .QN(n3134) );
  INVX0 U3175 ( .INP(n3135), .ZN(n3131) );
  XOR2X1 U3176 ( .IN1(n3136), .IN2(keyinput32), .Q(n3126) );
  NAND2X0 U3177 ( .IN1(n3137), .IN2(n3138), .QN(n3136) );
  XOR2X1 U3178 ( .IN1(n3139), .IN2(keyinput7), .Q(n3123) );
  NAND2X0 U3179 ( .IN1(N69), .IN2(N324), .QN(n3139) );
  XOR2X1 U3180 ( .IN1(n3140), .IN2(keyinput4), .Q(n3117) );
  NAND2X0 U3181 ( .IN1(N52), .IN2(N341), .QN(n3140) );
  INVX0 U3182 ( .INP(n3141), .ZN(n3103) );
  NAND2X0 U3183 ( .IN1(n3141), .IN2(n3142), .QN(N3211) );
  NAND3X0 U3184 ( .IN1(N375), .IN2(n3143), .IN3(N1), .QN(n3142) );
  AO21X1 U3185 ( .IN1(N1), .IN2(N375), .IN3(n3143), .Q(n3141) );
  AO21X1 U3186 ( .IN1(n3144), .IN2(n3145), .IN3(n3102), .Q(n3143) );
  NOR2X0 U3187 ( .IN1(n3145), .IN2(n3144), .QN(n3102) );
  NAND2X0 U3188 ( .IN1(n3107), .IN2(n3146), .QN(n3145) );
  NAND3X0 U3189 ( .IN1(N358), .IN2(n3147), .IN3(N18), .QN(n3146) );
  AO21X1 U3190 ( .IN1(N18), .IN2(N358), .IN3(n3147), .Q(n3107) );
  NAND2X0 U3191 ( .IN1(n3108), .IN2(n3148), .QN(n3147) );
  NAND3X0 U3192 ( .IN1(n3149), .IN2(n3150), .IN3(n3151), .QN(n3148) );
  AO21X1 U3193 ( .IN1(n3151), .IN2(n3150), .IN3(n3149), .Q(n3108) );
  NAND2X0 U3194 ( .IN1(n3114), .IN2(n3152), .QN(n3149) );
  NAND3X0 U3195 ( .IN1(N341), .IN2(n3153), .IN3(N35), .QN(n3152) );
  AO21X1 U3196 ( .IN1(N35), .IN2(N341), .IN3(n3153), .Q(n3114) );
  NAND2X0 U3197 ( .IN1(n3115), .IN2(n3154), .QN(n3153) );
  NAND3X0 U3198 ( .IN1(n3155), .IN2(n3156), .IN3(n3157), .QN(n3154) );
  AO21X1 U3199 ( .IN1(n3155), .IN2(n3156), .IN3(n3157), .Q(n3115) );
  NAND2X0 U3200 ( .IN1(n3120), .IN2(n3158), .QN(n3157) );
  NAND3X0 U3201 ( .IN1(N324), .IN2(n3159), .IN3(N52), .QN(n3158) );
  AO21X1 U3202 ( .IN1(N52), .IN2(N324), .IN3(n3159), .Q(n3120) );
  NAND2X0 U3203 ( .IN1(n3121), .IN2(n3160), .QN(n3159) );
  NAND3X0 U3204 ( .IN1(n3161), .IN2(n3162), .IN3(n3163), .QN(n3160) );
  AO21X1 U3205 ( .IN1(n3161), .IN2(n3162), .IN3(n3163), .Q(n3121) );
  NAND2X0 U3206 ( .IN1(n3138), .IN2(n3164), .QN(n3163) );
  NAND4X0 U3207 ( .IN1(n3165), .IN2(N69), .IN3(N307), .IN4(n3166), .QN(n3164)
         );
  AO22X1 U3208 ( .IN1(N69), .IN2(N307), .IN3(n3165), .IN4(n3166), .Q(n3138) );
  NAND2X0 U3209 ( .IN1(n3137), .IN2(n3167), .QN(n3166) );
  XOR2X1 U3210 ( .IN1(n3168), .IN2(keyinput27), .Q(n3165) );
  NAND2X0 U3211 ( .IN1(n3169), .IN2(n3137), .QN(n3168) );
  NAND2X0 U3212 ( .IN1(n3169), .IN2(n3167), .QN(n3137) );
  NAND3X0 U3213 ( .IN1(N273), .IN2(n3170), .IN3(N86), .QN(n3167) );
  AND2X1 U3214 ( .IN1(n3132), .IN2(n3171), .Q(n3169) );
  NAND3X0 U3215 ( .IN1(N290), .IN2(n3135), .IN3(N86), .QN(n3171) );
  AO21X1 U3216 ( .IN1(N86), .IN2(N290), .IN3(n3135), .Q(n3132) );
  NAND2X0 U3217 ( .IN1(N103), .IN2(N273), .QN(n3135) );
  INVX0 U3218 ( .INP(n3172), .ZN(n3162) );
  INVX0 U3219 ( .INP(n3173), .ZN(n3151) );
  XOR2X1 U3220 ( .IN1(n3174), .IN2(keyinput48), .Q(n3144) );
  NAND2X0 U3221 ( .IN1(n3175), .IN2(n3176), .QN(n3174) );
  INVX0 U3222 ( .INP(n3177), .ZN(n3176) );
  AO21X1 U3223 ( .IN1(n3178), .IN2(n3179), .IN3(n3177), .Q(N2877) );
  NOR2X0 U3224 ( .IN1(n3179), .IN2(n3178), .QN(n3177) );
  NAND2X0 U3225 ( .IN1(n3175), .IN2(n3180), .QN(n3179) );
  NAND3X0 U3226 ( .IN1(n3181), .IN2(n3182), .IN3(n3183), .QN(n3180) );
  AO21X1 U3227 ( .IN1(n3181), .IN2(n3182), .IN3(n3183), .Q(n3175) );
  AO21X1 U3228 ( .IN1(n3184), .IN2(n3185), .IN3(n3173), .Q(n3183) );
  NOR2X0 U3229 ( .IN1(n3185), .IN2(n3184), .QN(n3173) );
  NAND2X0 U3230 ( .IN1(n3150), .IN2(n3186), .QN(n3185) );
  NAND3X0 U3231 ( .IN1(n3187), .IN2(n3188), .IN3(n3189), .QN(n3186) );
  AO21X1 U3232 ( .IN1(n3187), .IN2(n3188), .IN3(n3189), .Q(n3150) );
  XOR2X1 U3233 ( .IN1(n3190), .IN2(keyinput37), .Q(n3189) );
  NAND2X0 U3234 ( .IN1(n3155), .IN2(n3191), .QN(n3190) );
  NAND3X0 U3235 ( .IN1(N324), .IN2(n3192), .IN3(N35), .QN(n3191) );
  AO21X1 U3236 ( .IN1(N35), .IN2(N324), .IN3(n3192), .Q(n3155) );
  NAND2X0 U3237 ( .IN1(n3156), .IN2(n3193), .QN(n3192) );
  NAND4X0 U3238 ( .IN1(n3194), .IN2(n3195), .IN3(n3196), .IN4(n3197), .QN(
        n3193) );
  AO22X1 U3239 ( .IN1(n3194), .IN2(n3196), .IN3(n3195), .IN4(n3197), .Q(n3156)
         );
  NAND2X0 U3240 ( .IN1(n3198), .IN2(n3161), .QN(n3196) );
  XNOR2X1 U3241 ( .IN1(n3199), .IN2(keyinput31), .Q(n3194) );
  NAND2X0 U3242 ( .IN1(n3161), .IN2(n3200), .QN(n3199) );
  NAND2X0 U3243 ( .IN1(n3198), .IN2(n3200), .QN(n3161) );
  NAND2X0 U3244 ( .IN1(N52), .IN2(N307), .QN(n3200) );
  AOI21X1 U3245 ( .IN1(n3201), .IN2(n3202), .IN3(n3172), .QN(n3198) );
  NOR2X0 U3246 ( .IN1(n3202), .IN2(n3201), .QN(n3172) );
  NAND2X0 U3247 ( .IN1(n3170), .IN2(n3203), .QN(n3202) );
  NAND3X0 U3248 ( .IN1(N69), .IN2(N290), .IN3(n3204), .QN(n3203) );
  AO21X1 U3249 ( .IN1(N69), .IN2(N290), .IN3(n3204), .Q(n3170) );
  XOR2X1 U3250 ( .IN1(n3205), .IN2(keyinput22), .Q(n3204) );
  NAND2X0 U3251 ( .IN1(N86), .IN2(N273), .QN(n3205) );
  XNOR2X1 U3252 ( .IN1(n3206), .IN2(keyinput2), .Q(n3184) );
  NAND2X0 U3253 ( .IN1(N18), .IN2(N341), .QN(n3206) );
  XNOR2X1 U3254 ( .IN1(n3207), .IN2(keyinput0), .Q(n3178) );
  NAND2X0 U3255 ( .IN1(N1), .IN2(N358), .QN(n3207) );
  NAND2X0 U3256 ( .IN1(n3181), .IN2(n3208), .QN(N2548) );
  NAND3X0 U3257 ( .IN1(N341), .IN2(n3209), .IN3(N1), .QN(n3208) );
  AO21X1 U3258 ( .IN1(N1), .IN2(N341), .IN3(n3209), .Q(n3181) );
  NAND2X0 U3259 ( .IN1(n3182), .IN2(n3210), .QN(n3209) );
  NAND3X0 U3260 ( .IN1(n3211), .IN2(n3212), .IN3(n3213), .QN(n3210) );
  AO21X1 U3261 ( .IN1(n3211), .IN2(n3212), .IN3(n3213), .Q(n3182) );
  NAND2X0 U3262 ( .IN1(n3187), .IN2(n3214), .QN(n3213) );
  NAND3X0 U3263 ( .IN1(N324), .IN2(n3215), .IN3(N18), .QN(n3214) );
  AO21X1 U3264 ( .IN1(N18), .IN2(N324), .IN3(n3215), .Q(n3187) );
  NAND2X0 U3265 ( .IN1(n3188), .IN2(n3216), .QN(n3215) );
  NAND3X0 U3266 ( .IN1(n3217), .IN2(n3218), .IN3(n3219), .QN(n3216) );
  AO21X1 U3267 ( .IN1(n3217), .IN2(n3218), .IN3(n3219), .Q(n3188) );
  NAND2X0 U3268 ( .IN1(n3195), .IN2(n3220), .QN(n3219) );
  NAND3X0 U3269 ( .IN1(N307), .IN2(n3221), .IN3(N35), .QN(n3220) );
  AO21X1 U3270 ( .IN1(N35), .IN2(N307), .IN3(n3221), .Q(n3195) );
  OAI21X1 U3271 ( .IN1(n3222), .IN2(n3201), .IN3(n3197), .QN(n3221) );
  AO21X1 U3272 ( .IN1(n3223), .IN2(n3224), .IN3(n3225), .Q(n3197) );
  AO21X1 U3273 ( .IN1(N52), .IN2(N290), .IN3(n3226), .Q(n3223) );
  INVX0 U3274 ( .INP(n3227), .ZN(n3226) );
  INVX0 U3275 ( .INP(n3224), .ZN(n3201) );
  NAND3X0 U3276 ( .IN1(N273), .IN2(n3227), .IN3(N69), .QN(n3224) );
  NAND3X0 U3277 ( .IN1(N273), .IN2(n3228), .IN3(N69), .QN(n3227) );
  NAND2X0 U3278 ( .IN1(N52), .IN2(N290), .QN(n3228) );
  NAND2X0 U3279 ( .IN1(n3211), .IN2(n3229), .QN(N2223) );
  NAND3X0 U3280 ( .IN1(N324), .IN2(n3230), .IN3(N1), .QN(n3229) );
  AO21X1 U3281 ( .IN1(N1), .IN2(N324), .IN3(n3230), .Q(n3211) );
  NAND2X0 U3282 ( .IN1(n3212), .IN2(n3231), .QN(n3230) );
  NAND3X0 U3283 ( .IN1(n3232), .IN2(n3233), .IN3(n3234), .QN(n3231) );
  AO21X1 U3284 ( .IN1(n3232), .IN2(n3233), .IN3(n3234), .Q(n3212) );
  XOR2X1 U3285 ( .IN1(n3235), .IN2(keyinput34), .Q(n3234) );
  NAND2X0 U3286 ( .IN1(n3217), .IN2(n3236), .QN(n3235) );
  NAND3X0 U3287 ( .IN1(N307), .IN2(n3237), .IN3(N18), .QN(n3236) );
  AO21X1 U3288 ( .IN1(N18), .IN2(N307), .IN3(n3237), .Q(n3217) );
  OAI21X1 U3289 ( .IN1(n3238), .IN2(n3225), .IN3(n3218), .QN(n3237) );
  AO21X1 U3290 ( .IN1(n3239), .IN2(n3222), .IN3(n3240), .Q(n3218) );
  INVX0 U3291 ( .INP(n3238), .ZN(n3240) );
  AO21X1 U3292 ( .IN1(N35), .IN2(N290), .IN3(n3241), .Q(n3239) );
  INVX0 U3293 ( .INP(n3242), .ZN(n3241) );
  INVX0 U3294 ( .INP(n3222), .ZN(n3225) );
  NAND3X0 U3295 ( .IN1(N273), .IN2(n3242), .IN3(N52), .QN(n3222) );
  NAND3X0 U3296 ( .IN1(N273), .IN2(n3243), .IN3(N52), .QN(n3242) );
  NAND2X0 U3297 ( .IN1(N35), .IN2(N290), .QN(n3243) );
  INVX0 U3298 ( .INP(n3244), .ZN(n3233) );
  NAND2X0 U3299 ( .IN1(n3232), .IN2(n3245), .QN(N1901) );
  NAND3X0 U3300 ( .IN1(N307), .IN2(n3246), .IN3(N1), .QN(n3245) );
  AO21X1 U3301 ( .IN1(N1), .IN2(N307), .IN3(n3246), .Q(n3232) );
  AO21X1 U3302 ( .IN1(n3247), .IN2(n3248), .IN3(n3244), .Q(n3246) );
  NOR2X0 U3303 ( .IN1(n3248), .IN2(n3247), .QN(n3244) );
  XOR2X1 U3304 ( .IN1(n3249), .IN2(keyinput24), .Q(n3248) );
  AND2X1 U3305 ( .IN1(n3250), .IN2(n3238), .Q(n3247) );
  NAND3X0 U3306 ( .IN1(N273), .IN2(n3251), .IN3(N35), .QN(n3238) );
  AO21X1 U3307 ( .IN1(N18), .IN2(N290), .IN3(n3252), .Q(n3250) );
  INVX0 U3308 ( .INP(n3251), .ZN(n3252) );
  NAND3X0 U3309 ( .IN1(N273), .IN2(n3253), .IN3(N35), .QN(n3251) );
  NAND2X0 U3310 ( .IN1(N18), .IN2(N290), .QN(n3253) );
  OA21X1 U3311 ( .IN1(n3254), .IN2(n3255), .IN3(n3249), .Q(N1581) );
  NAND3X0 U3312 ( .IN1(N273), .IN2(n3256), .IN3(N18), .QN(n3249) );
  INVX0 U3313 ( .INP(n3256), .ZN(n3255) );
  NAND3X0 U3314 ( .IN1(N273), .IN2(n3257), .IN3(N18), .QN(n3256) );
  NAND2X0 U3315 ( .IN1(N1), .IN2(N290), .QN(n3257) );
  NOR2X0 U3316 ( .IN1(n2925), .IN2(n2601), .QN(n3254) );
  INVX0 U3317 ( .INP(N1), .ZN(n2601) );
  INVX0 U3318 ( .INP(N290), .ZN(n2925) );
endmodule

