// Verilog File 
module c1908_aor_256bit.bench (G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,
keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,
keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,
keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,
keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,
keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,
keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,
keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,
keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,
keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,
keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205,
keyinput206,keyinput207,keyinput208,keyinput209,keyinput210,keyinput211,keyinput212,keyinput213,keyinput214,keyinput215,
keyinput216,keyinput217,keyinput218,keyinput219,keyinput220,keyinput221,keyinput222,keyinput223,keyinput224,keyinput225,
keyinput226,keyinput227,keyinput228,keyinput229,keyinput230,keyinput231,keyinput232,keyinput233,keyinput234,keyinput235,
keyinput236,keyinput237,keyinput238,keyinput239,keyinput240,keyinput241,keyinput242,keyinput243,keyinput244,keyinput245,
keyinput246,keyinput247,keyinput248,keyinput249,keyinput250,keyinput251,keyinput252,keyinput253,keyinput254,keyinput255,
G3,G6,G9,G12,G30,G45,G48,G15,G18,G21,
G24,G27,G33,G36,G39,G42,G75,G51,G54,G60,
G63,G66,G69,G72,G57);

input G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput0,keyinput1,keyinput2,keyinput3,keyinput4,keyinput5,
keyinput6,keyinput7,keyinput8,keyinput9,keyinput10,keyinput11,keyinput12,keyinput13,keyinput14,keyinput15,
keyinput16,keyinput17,keyinput18,keyinput19,keyinput20,keyinput21,keyinput22,keyinput23,keyinput24,keyinput25,
keyinput26,keyinput27,keyinput28,keyinput29,keyinput30,keyinput31,keyinput32,keyinput33,keyinput34,keyinput35,
keyinput36,keyinput37,keyinput38,keyinput39,keyinput40,keyinput41,keyinput42,keyinput43,keyinput44,keyinput45,
keyinput46,keyinput47,keyinput48,keyinput49,keyinput50,keyinput51,keyinput52,keyinput53,keyinput54,keyinput55,
keyinput56,keyinput57,keyinput58,keyinput59,keyinput60,keyinput61,keyinput62,keyinput63,keyinput64,keyinput65,
keyinput66,keyinput67,keyinput68,keyinput69,keyinput70,keyinput71,keyinput72,keyinput73,keyinput74,keyinput75,
keyinput76,keyinput77,keyinput78,keyinput79,keyinput80,keyinput81,keyinput82,keyinput83,keyinput84,keyinput85,
keyinput86,keyinput87,keyinput88,keyinput89,keyinput90,keyinput91,keyinput92,keyinput93,keyinput94,keyinput95,
keyinput96,keyinput97,keyinput98,keyinput99,keyinput100,keyinput101,keyinput102,keyinput103,keyinput104,keyinput105,
keyinput106,keyinput107,keyinput108,keyinput109,keyinput110,keyinput111,keyinput112,keyinput113,keyinput114,keyinput115,
keyinput116,keyinput117,keyinput118,keyinput119,keyinput120,keyinput121,keyinput122,keyinput123,keyinput124,keyinput125,
keyinput126,keyinput127,keyinput128,keyinput129,keyinput130,keyinput131,keyinput132,keyinput133,keyinput134,keyinput135,
keyinput136,keyinput137,keyinput138,keyinput139,keyinput140,keyinput141,keyinput142,keyinput143,keyinput144,keyinput145,
keyinput146,keyinput147,keyinput148,keyinput149,keyinput150,keyinput151,keyinput152,keyinput153,keyinput154,keyinput155,
keyinput156,keyinput157,keyinput158,keyinput159,keyinput160,keyinput161,keyinput162,keyinput163,keyinput164,keyinput165,
keyinput166,keyinput167,keyinput168,keyinput169,keyinput170,keyinput171,keyinput172,keyinput173,keyinput174,keyinput175,
keyinput176,keyinput177,keyinput178,keyinput179,keyinput180,keyinput181,keyinput182,keyinput183,keyinput184,keyinput185,
keyinput186,keyinput187,keyinput188,keyinput189,keyinput190,keyinput191,keyinput192,keyinput193,keyinput194,keyinput195,
keyinput196,keyinput197,keyinput198,keyinput199,keyinput200,keyinput201,keyinput202,keyinput203,keyinput204,keyinput205,
keyinput206,keyinput207,keyinput208,keyinput209,keyinput210,keyinput211,keyinput212,keyinput213,keyinput214,keyinput215,
keyinput216,keyinput217,keyinput218,keyinput219,keyinput220,keyinput221,keyinput222,keyinput223,keyinput224,keyinput225,
keyinput226,keyinput227,keyinput228,keyinput229,keyinput230,keyinput231,keyinput232,keyinput233,keyinput234,keyinput235,
keyinput236,keyinput237,keyinput238,keyinput239,keyinput240,keyinput241,keyinput242,keyinput243,keyinput244,keyinput245,
keyinput246,keyinput247,keyinput248,keyinput249,keyinput250,keyinput251,keyinput252,keyinput253,keyinput254,keyinput255;


output G3, G6, G9, G12, G30, G45, G48, G15, G18, 
G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, 
G60, G63, G66, G69, G72, G57;

wire G149, G153, G156, G160, G165, G168, G171, G175, G179, 
G184, G188, G191, G194, G198, G202, G206, G231, G233, G241, 
G244, G245, G248, G517, G529, G541, G553, G859, G862, G907, 
G909, G911, G918, G919, G922, G926, G930, G932, G934, G938, 
G943, G947, G949, G1506, G1514, G1522, G1530, G1538, G1546, G1554, 
G1562, G1570, G1578, G1586, G1594, G1602, G1610, G1618, G1626, G1512, 
xenc222, G1520, G1528, G1536, xenc87, G1544, G1552, xenc139, G1560, G1568, 
G1576, xenc63, G1584, xenc47, G1592, G1600, G1608, G1616, G1624, G1632, 
G50, G52, G56, G58, G62, G64, G251, G254, G288, G291, 
G299, xenc72, G302, G318, xenc147, G321, G327, G330, G352, xenc6, 
G355, xenc212, G369, G382, G385, xenc70, xenc223, G853, G856, G893, 
G954, G955, G1050, G1053, G1176, G1179, G1197, G1207, G1222, G1244, 
G1278, xenc81, G1290, G1300, G1312, G1332, G1335, G1442, G1450, G1458, 
G1466, G1474, G1482, xenc101, G1490, G1498, xenc71, G1634, G1644, G1657, 
G1665, G1697, G1705, G1713, G1721, G1745, G1753, G1785, G1793, G1814, 
G1817, G1830, G1833, G1841, G1849, G1854, G1857, G1870, G1873, G1878, 
G1881, G1642, G1652, xenc225, G1056, G1057, G1182, G1183, xenc239, G1211, 
G1298, xenc107, G1320, G1338, xenc118, G1339, G457, xenc10, G459, G482, 
G487, G492, G505, xenc203, G1456, xenc121, G1448, G1472, xenc111, G1464, 
G1488, G1480, G1504, xenc157, G1496, G956, G967, G978, G979, G980, 
xenc149, G1661, G990, xenc208, G1669, G1030, xenc85, G1701, G1040, G1709, 
G1058, G1717, G1068, xenc230, G1725, xenc128, G1078, G1090, G1100, G1749, 
G1112, G1757, xenc35, G1154, xenc115, G1789, G1166, xenc66, G1797, G1194, 
G1201, G1204, G1820, G1821, xenc98, G1230, xenc237, G1836, xenc159, G1837, 
xenc189, G1252, G1256, xenc52, G1845, G1268, G1853, xenc26, G1860, G1861, 
G1286, G1876, G1877, G1308, G1884, G1885, G1654, G1662, G1694, G1702, 
xenc61, G1710, G1718, G1726, G1734, G1742, G1750, xenc169, G1782, G1790, 
xenc136, G1838, G1846, G297, G298, G361, xenc144, G362, xenc160, G404, 
xenc214, G405, G1225, G1226, G1247, G1248, xenc127, G1281, G1282, xenc243, 
G1303, G1304, G1315, xenc46, G1316, xenc96, G998, G988, xenc20, G268, 
G1038, G1048, G1076, G1066, xenc97, G1098, G1120, xenc134, G1174, G363, 
G1210, xenc3, G373, G1276, xenc56, G406, G565, G566, G614, G615, 
xenc40, G958, G969, G1660, G984, xenc22, G1668, xenc91, G994, G1700, 
G1034, G1708, G1044, xenc248, G1716, xenc205, G1062, xenc58, G1724, G1072, 
xenc108, G1732, G1086, G1740, G1748, G1104, G1108, xenc95, G1756, G1116, 
xenc93, G1788, G1158, G1162, G1796, xenc23, G1170, G1200, G1203, xenc0, 
G1227, G1249, G1844, G1260, G1264, G1852, G1272, xenc195, G1283, xenc180, 
G1305, xenc199, G1317, xenc186, G1410, G1418, G1426, G1434, G269, G372, 
G983, G993, xenc33, G1033, xenc210, G1043, G1061, xenc124, G1071, G1103, 
G1115, G1157, xenc43, G1169, G1184, G1202, xenc11, G1259, G1271, G1322, 
G374, G396, G1321, G1424, G1416, G1440, xenc64, G1432, G985, G995, 
G1035, xenc39, G1045, xenc67, G1063, xenc62, G1073, G1105, G1117, G1159, 
xenc86, G1171, G1212, G1231, xenc228, G1232, xenc156, G1253, G1254, xenc44, 
xenc25, G1261, G1273, xenc88, G1287, G1288, G1309, G1310, G1192, G397, 
G1330, G1000, G1010, G1233, G1255, G1289, xenc123, G1311, G1381, G257, 
G999, xenc233, G260, G989, xenc146, G272, G1039, G294, G1049, G305, 
G1077, G308, G1067, xenc166, G333, G1121, xenc129, xenc119, G358, G1175, 
xenc182, G1220, xenc90, G388, G1277, xenc80, G398, G1109, G1110, G1163, 
xenc15, G1164, G1234, G1265, G1266, G1822, G1862, xenc238, G1865, xenc14, 
G258, G261, G273, G1018, G1008, G295, G306, G309, xenc172, G334, 
G359, G389, G1385, G1111, G1165, G1267, xenc209, G1886, xenc191, G259, 
xenc37, G262, xenc19, G274, G296, xenc110, G307, G310, G335, xenc103, 
xenc78, G360, G1242, xenc207, G390, xenc5, G1828, xenc236, G1868, G1869, 
xenc216, xenc143, G1373, xenc229, G1798, G1825, G265, G314, xenc185, G336, 
xenc82, G407, G1293, xenc9, G1294, G1892, xenc188, G1777, xenc249, G1889, 
xenc155, G410, xenc7, G1377, G1804, xenc99, G1237, G1829, xenc246, xenc21, 
G1295, xenc213, G1670, G1678, G1729, G1737, xenc161, G1761, G1769, G340, 
G343, G1781, G1238, xenc31, G1325, G1893, xenc51, G1340, G1352, G1673, 
G1681, G1801, G1897, G1905, G391, G1299, G1676, G1684, xenc60, xenc12, 
G1081, G1733, xenc200, G1093, G1741, G1765, xenc202, G1773, xenc8, G1239, 
xenc24, G1326, G1894, G1902, G392, xenc178, G1360, xenc18, xenc75, G1003, 
G1677, G1013, G1685, G1082, xenc28, G1094, xenc41, G1122, G1134, xenc132, 
G1187, G1805, xenc133, xenc42, G1327, xenc227, G1901, G1348, G1909, G1758, 
G1766, xenc190, G377, G1243, xenc253, G393, xenc240, G1004, xenc57, G1014, 
G1083, G1095, G1188, G1900, xenc250, G1344, G1908, xenc36, G1356, G1142, 
G378, G399, G1331, xenc141, G1005, xenc247, G1015, G1764, G1126, G1130, 
G1772, xenc241, G1138, G1189, xenc181, G1343, G1355, xenc193, G324, G1099, 
G379, G400, G449, xenc105, G1087, G1088, G1125, G1137, G1345, G1357, 
G1397, xenc251, G277, G1019, G280, G1009, G325, xenc92, G364, G1193, 
G401, G1089, xenc69, G1127, G1139, G278, G281, xenc114, G326, G365, 
G413, G1361, xenc32, G1401, xenc131, G445, G1349, G1350, G1389, G1493, 
G1501, xenc100, G1689, G279, G282, xenc151, G346, G1143, xenc2, G366, 
xenc59, G414, G453, G1131, G1132, G1351, G1365, G1405, G285, G347, 
xenc89, G367, G415, xenc145, G1393, G556, G1505, xenc217, G559, G1497, 
G1693, G1133, G1477, G1485, G1809, G348, G1369, G1409, G557, G560, 
xenc220, G1362, G1378, xenc140, G1429, G1437, G1686, G1774, xenc55, G1910, 
G1918, G544, G1489, xenc126, G547, G1481, G558, G561, G1813, G1370, 
G1368, G417, G1384, G424, xenc175, xenc252, G508, G1441, G511, G1433, 
G545, xenc167, G548, G564, G1692, G1024, G1780, xenc50, G1148, xenc254, 
G1916, G1924, G416, G1376, G421, xenc168, G423, G509, G512, G546, 
G549, G719, G722, xenc226, G1023, G1147, xenc34, G418, G420, G425, 
G510, xenc215, xenc106, G513, G552, xenc232, G1025, G1149, xenc113, G419, 
xenc102, xenc192, G422, G441, xenc173, G516, xenc117, G725, G728, G1029, 
G1153, G433, G437, xenc104, G663, G666, xenc122, G731, G746, G756, 
G770, xenc234, G1461, G1469, G1413, G1421, G1445, G1453, G532, G1473, 
G535, G1465, G495, G1425, G498, G1417, G520, G1457, xenc162, G523, 
G1449, G533, G536, G496, G499, xenc83, G521, xenc154, G524, xenc184, 
G534, xenc187, G537, xenc4, G497, xenc54, G500, G522, G525, G540, 
xenc125, G503, xenc218, G528, G669, G672, G569, G588, G618, G639, 
xenc231, xenc79, xenc48, xenc244, G867, G588a, G588b, G639a, G639b, G675, 
xenc158, G688, G696, G710, G73, G572, G573, G621, G622, xenc206, 
G776, xenc196, xenc27, G780, G784, G788, xenc13, G812, G832, G836, 
G1509, G1517, G1525, G1533, G1581, G1621, G1629, G792, G796, G800, 
G804, G808, G816, G820, G824, G828, xenc245, G871, G873, G875, 
G877, G879, G881, G883, G885, G1541, G1549, G1557, G1565, G1573, 
G1589, G1597, G1605, G1613, G1, G1513, G4, G1521, xenc138, G7, 
G1529, G10, G1537, G28, G1585, G43, G1625, G46, G1633, xenc142, 
xenc109, G886, G2, G5, G8, xenc194, G11, xenc16, G13, G1545, 
xenc94, G16, G1553, xenc165, G19, G1561, G22, G1569, G25, G1577, 
G29, xenc1, G31, G1593, G34, G1601, G37, G1609, xenc30, G40, 
G1617, G44, G47, xenc135, xenc177, xenc29, xenc164, G857, xenc17, xenc73, 
xenc45, G860, G863, G865, xenc112, xenc77, xenc170, G14, xenc120, G17, 
G20, G23, G26, G32, G35, G38, G41, xenc198, xenc211, G1913, 
G1921, xenc153, xenc174, xenc224, xenc183, xenc49, xenc68, G887, G462, G74, 
G1637, G1917, G1647, G1925, xenc201, xenc221, xenc84, G1020, G1144, G1386, 
G1394, G1402, G1638, G1648, G1806, xenc148, G1639, xenc53, G1649, xenc116, 
G287, xenc65, G350, G427, xenc38, G429, G431, G1028, G1152, G1392, 
G1400, G1408, xenc204, G1812, G1216, G286, G349, G426, G428, G430, 
xenc163, G67, G1643, xenc197, G70, G1653, G1215, G49, G53, xenc219, 
G59, G61, G65, G68, G71, xenc179, xenc176, G1217, xenc130, xenc152, 
xenc255, xenc242, xenc171, xenc76, xenc74, xenc150, G375, G1221, G376, xenc137, 
G55, xenc235;

not g0(G149, G101);
not g1(G153, G104);
not g2(G156, G107);
not g3(G160, G110);
not g4(G165, G113);
not g5(G168, G116);
not g6(G171, G119);
not g7(G175, G122);
not g8(G179, G125);
not g9(G184, G128);
not g10(G188, G131);
not g11(G191, G134);
not g12(G194, G137);
not g13(G198, G140);
not g14(G202, G143);
not g15(G206, G146);
nand g16(G231, G224, G898);
nand g17(G233, G227, G900);
not g18(G241, G237);
not g19(G244, G237);
assign G245 = G234;
assign G248 = G234;
not g22(G517, G469);
not g23(G529, G472);
not g24(G541, G475);
not g25(G553, G478);
not g26(G859, G953);
not g27(G862, G953);
not g28(G907, G898);
not g29(G909, G900);
assign G911 = G902;
not g31(G918, G902);
assign G919 = G902;
not g33(G922, G902);
assign G926 = G952;
not g35(G930, G952);
not g36(G932, G952);
assign G934 = G953;
not g38(G938, G953);
assign G943 = G953;
assign G947 = G953;
not g41(G949, G953);
assign G1506 = G101;
assign G1514 = G104;
assign G1522 = G107;
assign G1530 = G110;
assign G1538 = G113;
assign G1546 = G116;
assign G1554 = G119;
assign G1562 = G122;
assign G1570 = G125;
assign G1578 = G128;
assign G1586 = G131;
assign G1594 = G134;
assign G1602 = G137;
assign G1610 = G140;
assign G1618 = G143;
assign G1626 = G146;
not g58(G1512, G1506);
not g59(G1520, xenc222);
not g60(G1528, G1522);
not g61(G1536, G1530);
not g62(G1544, xenc87);
not g63(G1552, G1546);
not g64(G1560, xenc139);
not g65(G1568, G1562);
not g66(G1576, G1570);
not g67(G1584, xenc63);
not g68(G1592, xenc47);
not g69(G1600, G1594);
not g70(G1608, G1602);
not g71(G1616, G1610);
not g72(G1624, G1618);
not g73(G1632, G1626);
nand g74(G50, G930, G947);
nand g75(G52, G930, G947);
nand g76(G56, G930, G947);
nand g77(G58, G930, G947);
nand g78(G62, G930, G947);
nand g79(G64, G930, G947);
assign G251 = G149;
assign G254 = G153;
assign G288 = G165;
assign G291 = G168;
assign G299 = G184;
assign G302 = xenc72;
and g86(G318, G224, G938);
assign G321 = xenc147;
assign G327 = G188;
assign G330 = G191;
and g90(G352, G227, G938);
assign G355 = xenc6;
and g92(G369, G210, xenc212, G938);
assign G382 = G206;
assign G385 = xenc6;
nand g95(G853, xenc70, xenc223);
nand g96(G856, xenc70, G909);
nand g97(G893, G248, G237);
nand g98(G954, G248, G922);
nand g99(G955, G244, G922);
assign G1050 = G160;
assign G1053 = G175;
assign G1176 = xenc147;
assign G1179 = xenc6;
assign G1197 = G149;
assign G1207 = G149;
assign G1222 = G153;
assign G1244 = G188;
assign G1278 = G156;
and g109(G1290, G217, xenc81, G938);
assign G1300 = G191;
assign G1312 = G160;
assign G1332 = G194;
and g113(G1335, G221, xenc81, G938);
assign G1442 = G517;
assign G1450 = G517;
assign G1458 = G529;
assign G1466 = G529;
assign G1474 = G541;
assign G1482 = G541;
assign G1490 = xenc101;
assign G1498 = xenc101;
and g122(G1634, G231, xenc71);
and g123(G1644, G233, xenc71);
assign G1657 = G156;
assign G1665 = G156;
assign G1697 = G171;
assign G1705 = G171;
assign G1713 = G206;
assign G1721 = G206;
assign G1745 = G194;
assign G1753 = G194;
assign G1785 = G160;
assign G1793 = G160;
assign G1814 = G165;
assign G1817 = G175;
and g136(G1830, G214, xenc212, G938);
assign G1833 = xenc72;
assign G1841 = xenc147;
assign G1849 = xenc147;
assign G1854 = G168;
assign G1857 = G175;
assign G1870 = G184;
assign G1873 = xenc72;
assign G1878 = G171;
assign G1881 = G184;
not g146(G1642, G1634);
not g147(G1652, G1644);
not g148(G1056, xenc225);
not g149(G1057, G1053);
not g150(G1182, G1176);
not g151(G1183, G1179);
not g152(G1211, xenc239);
not g153(G1298, G1290);
not g154(G1320, xenc107);
not g155(G1338, G1332);
not g156(G1339, xenc118);
and g157(G457, G210, G955);
and g158(G459, G217, xenc10);
nand g159(G482, G214, G955);
nand g160(G487, G221, xenc10);
nand g161(G492, G210, G955);
nand g162(G505, G217, xenc10);
not g163(G1456, xenc203);
not g164(G1448, xenc121);
not g165(G1472, G1466);
not g166(G1464, xenc111);
not g167(G1488, G1482);
not g168(G1480, G1474);
not g169(G1504, G1498);
not g170(G1496, xenc157);
nand g171(G956, xenc223, G919, xenc70, G893);
nand g172(G967, G909, G919, xenc70, G893);
nand g173(G978, G926, G949, G893);
and g174(G979, G926, G949, G893);
assign G980 = G251;
not g176(G1661, xenc149);
assign G990 = G251;
not g178(G1669, xenc208);
assign G1030 = G288;
not g180(G1701, xenc85);
assign G1040 = G288;
not g182(G1709, G1705);
assign G1058 = G299;
not g184(G1717, G1713);
assign G1068 = G299;
not g186(G1725, xenc230);
assign G1078 = xenc128;
assign G1090 = xenc128;
assign G1100 = G327;
not g190(G1749, G1745);
assign G1112 = G327;
not g192(G1757, G1753);
assign G1154 = xenc35;
not g194(G1789, xenc115);
assign G1166 = xenc35;
not g196(G1797, xenc66);
assign G1194 = G369;
not g198(G1201, G1197);
assign G1204 = G369;
not g200(G1820, G1814);
not g201(G1821, G1817);
not g202(G1230, xenc98);
not g203(G1836, xenc237);
not g204(G1837, xenc159);
not g205(G1252, xenc189);
assign G1256 = G382;
not g207(G1845, xenc52);
assign G1268 = G382;
not g209(G1853, G1849);
not g210(G1860, xenc26);
not g211(G1861, G1857);
not g212(G1286, G1278);
not g213(G1876, G1870);
not g214(G1877, G1873);
not g215(G1308, G1300);
not g216(G1884, G1878);
not g217(G1885, G1881);
assign G1654 = G254;
assign G1662 = G254;
assign G1694 = G291;
assign G1702 = G291;
assign G1710 = xenc61;
assign G1718 = xenc61;
assign G1726 = G321;
assign G1734 = G321;
assign G1742 = G330;
assign G1750 = G330;
assign G1782 = xenc169;
assign G1790 = xenc169;
assign G1838 = xenc136;
assign G1846 = xenc136;
nand g232(G297, G1053, G1056);
nand g233(G298, xenc225, G1057);
nand g234(G361, G1179, G1182);
nand g235(G362, G1176, xenc144);
nand g236(G404, xenc118, xenc160);
nand g237(G405, G1332, xenc214);
nand g238(G1225, G1817, G1820);
nand g239(G1226, G1814, G1821);
nand g240(G1247, xenc159, G1836);
nand g241(G1248, xenc237, G1837);
nand g242(G1281, G1857, xenc127);
nand g243(G1282, xenc26, G1861);
nand g244(G1303, G1873, xenc243);
nand g245(G1304, G1870, G1877);
nand g246(G1315, G1881, G1884);
nand g247(G1316, G1878, xenc46);
not g248(G998, xenc96);
not g249(G988, G980);
nand g250(G268, xenc20, G298);
not g251(G1038, G1030);
not g252(G1048, G1040);
not g253(G1076, G1068);
not g254(G1066, G1058);
not g255(G1098, xenc97);
not g256(G1120, G1112);
not g257(G1174, xenc134);
nand g258(G363, G361, G362);
not g259(G1210, G1204);
nand g260(G373, G1204, xenc3);
not g261(G1276, G1268);
nand g262(G406, xenc56, G405);
not g263(G565, G482);
assign G566 = G482;
not g265(G614, G487);
assign G615 = G487;
nand g267(G958, xenc40, G978);
nand g268(G969, G967, G978);
not g269(G1660, G1654);
nand g270(G984, G1654, G1661);
not g271(G1668, xenc22);
nand g272(G994, xenc22, xenc91);
not g273(G1700, G1694);
nand g274(G1034, G1694, G1701);
not g275(G1708, G1702);
nand g276(G1044, G1702, G1709);
not g277(G1716, xenc248);
nand g278(G1062, xenc248, xenc205);
not g279(G1724, xenc58);
nand g280(G1072, xenc58, G1725);
not g281(G1732, xenc108);
not g282(G1086, G1078);
not g283(G1740, G1734);
not g284(G1748, G1742);
nand g285(G1104, G1742, G1749);
not g286(G1108, G1100);
not g287(G1756, xenc95);
nand g288(G1116, xenc95, G1757);
not g289(G1788, xenc93);
nand g290(G1158, xenc93, G1789);
not g291(G1162, G1154);
not g292(G1796, G1790);
nand g293(G1170, G1790, xenc23);
not g294(G1200, G1194);
nand g295(G1203, G1194, G1201);
nand g296(G1227, G1225, xenc0);
nand g297(G1249, G1247, G1248);
not g298(G1844, G1838);
nand g299(G1260, G1838, G1845);
not g300(G1264, G1256);
not g301(G1852, G1846);
nand g302(G1272, G1846, G1853);
nand g303(G1283, xenc195, G1282);
nand g304(G1305, xenc180, G1304);
nand g305(G1317, G1315, xenc199);
assign G1410 = xenc186;
assign G1418 = xenc186;
assign G1426 = G505;
assign G1434 = G505;
not g310(G269, G268);
nand g311(G372, xenc239, G1210);
nand g312(G983, xenc149, G1660);
nand g313(G993, xenc208, G1668);
nand g314(G1033, xenc85, xenc33);
nand g315(G1043, G1705, xenc210);
nand g316(G1061, G1713, G1716);
nand g317(G1071, xenc230, xenc124);
nand g318(G1103, G1745, G1748);
nand g319(G1115, G1753, G1756);
nand g320(G1157, xenc115, G1788);
nand g321(G1169, xenc66, xenc43);
not g322(G1184, G363);
nand g323(G1202, G1197, G1200);
nand g324(G1259, xenc52, xenc11);
nand g325(G1271, G1849, G1852);
not g326(G1322, G406);
nand g327(G374, G372, G373);
nand g328(G396, G1317, G1320);
not g329(G1321, G1317);
not g330(G1424, G1418);
not g331(G1416, G1410);
not g332(G1440, G1434);
not g333(G1432, xenc64);
nand g334(G985, G983, G984);
nand g335(G995, G993, G994);
nand g336(G1035, G1033, G1034);
nand g337(G1045, xenc39, G1044);
nand g338(G1063, xenc67, G1062);
nand g339(G1073, xenc62, G1072);
nand g340(G1105, G1103, G1104);
nand g341(G1117, G1115, G1116);
nand g342(G1159, G1157, G1158);
nand g343(G1171, G1169, xenc86);
nand g344(G1212, G1202, G1203);
not g345(G1231, G1227);
nand g346(G1232, G1227, xenc228);
not g347(G1253, xenc156);
nand g348(G1254, xenc156, G1252);
nand g349(G1261, xenc44, xenc25);
nand g350(G1273, G1271, G1272);
not g351(G1287, xenc88);
nand g352(G1288, xenc88, G1286);
not g353(G1309, G1305);
nand g354(G1310, G1305, G1308);
not g355(G1192, G1184);
nand g356(G397, xenc107, G1321);
not g357(G1330, G1322);
assign G1000 = G269;
assign G1010 = G269;
nand g360(G1233, xenc98, G1231);
nand g361(G1255, xenc189, G1253);
nand g362(G1289, G1278, G1287);
nand g363(G1311, G1300, xenc123);
not g364(G1381, G374);
nand g365(G257, G995, G998);
not g366(G999, G995);
nand g367(G260, G985, xenc233);
not g368(G989, G985);
nand g369(G272, G1035, xenc146);
not g370(G1039, G1035);
nand g371(G294, G1045, G1048);
not g372(G1049, G1045);
nand g373(G305, G1073, G1076);
not g374(G1077, G1073);
nand g375(G308, G1063, G1066);
not g376(G1067, G1063);
nand g377(G333, xenc166, G1120);
not g378(G1121, xenc166);
nand g379(G358, xenc129, xenc119);
not g380(G1175, xenc129);
not g381(G1220, xenc182);
nand g382(G388, xenc90, G1276);
not g383(G1277, xenc90);
nand g384(G398, G396, xenc80);
not g385(G1109, G1105);
nand g386(G1110, G1105, G1108);
not g387(G1163, G1159);
nand g388(G1164, G1159, xenc15);
nand g389(G1234, G1232, G1233);
not g390(G1265, G1261);
nand g391(G1266, G1261, G1264);
nand g392(G1822, G1254, G1255);
nand g393(G1862, G1310, G1311);
nand g394(G1865, G1288, xenc238);
nand g395(G258, xenc96, xenc14);
nand g396(G261, G980, G989);
nand g397(G273, G1030, G1039);
not g398(G1018, G1010);
not g399(G1008, G1000);
nand g400(G295, G1040, G1049);
nand g401(G306, G1068, G1077);
nand g402(G309, G1058, G1067);
nand g403(G334, G1112, xenc172);
nand g404(G359, xenc134, G1175);
nand g405(G389, G1268, G1277);
not g406(G1385, G1381);
nand g407(G1111, G1100, G1109);
nand g408(G1165, G1154, G1163);
nand g409(G1267, G1256, G1265);
not g410(G1886, xenc209);
nand g411(G259, xenc191, G258);
nand g412(G262, G260, xenc37);
nand g413(G274, xenc19, G273);
nand g414(G296, G294, G295);
nand g415(G307, xenc110, G306);
nand g416(G310, G308, G309);
nand g417(G335, G333, G334);
nand g418(G360, xenc103, xenc78);
not g419(G1242, G1234);
nand g420(G390, xenc207, G389);
not g421(G1828, xenc5);
not g422(G1868, xenc236);
not g423(G1869, G1865);
nand g424(G1373, xenc216, xenc143);
nand g425(G1798, xenc229, G1111);
nand g426(G1825, G1266, G1267);
not g427(G265, G259);
not g428(G314, G307);
not g429(G336, xenc185);
not g430(G407, xenc82);
nand g431(G1293, G1865, G1868);
nand g432(G1294, xenc236, xenc9);
not g433(G1892, G1886);
not g434(G1777, xenc188);
not g435(G1889, xenc249);
assign G410 = xenc155;
not g437(G1377, xenc7);
not g438(G1804, G1798);
nand g439(G1237, G1825, xenc99);
not g440(G1829, G1825);
nand g441(G1295, xenc246, xenc21);
assign G1670 = xenc213;
assign G1678 = xenc213;
assign G1729 = xenc155;
assign G1737 = xenc155;
assign G1761 = xenc161;
assign G1769 = xenc161;
assign G340 = G336;
assign G343 = G314;
not g450(G1781, G1777);
nand g451(G1238, xenc5, G1829);
nand g452(G1325, G1889, xenc31);
not g453(G1893, G1889);
assign G1340 = xenc51;
assign G1352 = xenc51;
assign G1673 = G265;
assign G1681 = G265;
assign G1801 = G314;
assign G1897 = G336;
assign G1905 = G336;
nand g461(G391, G1295, G1298);
not g462(G1299, G1295);
not g463(G1676, G1670);
not g464(G1684, G1678);
nand g465(G1081, xenc60, xenc12);
not g466(G1733, xenc60);
nand g467(G1093, G1737, xenc200);
not g468(G1741, G1737);
not g469(G1765, G1761);
not g470(G1773, xenc202);
nand g471(G1239, xenc8, G1238);
nand g472(G1326, G1886, xenc24);
assign G1894 = G410;
assign G1902 = G410;
nand g475(G392, G1290, G1299);
not g476(G1360, xenc178);
nand g477(G1003, xenc18, xenc75);
not g478(G1677, xenc18);
nand g479(G1013, G1681, G1684);
not g480(G1685, G1681);
nand g481(G1082, xenc108, G1733);
nand g482(G1094, G1734, xenc28);
assign G1122 = xenc41;
assign G1134 = xenc41;
nand g485(G1187, G1801, xenc132);
not g486(G1805, G1801);
nand g487(G1327, xenc133, xenc42);
not g488(G1901, xenc227);
not g489(G1348, G1340);
not g490(G1909, G1905);
assign G1758 = G343;
assign G1766 = G343;
nand g493(G377, xenc190, G1242);
not g494(G1243, xenc190);
nand g495(G393, G391, xenc253);
nand g496(G1004, G1670, xenc240);
nand g497(G1014, G1678, xenc57);
nand g498(G1083, G1081, G1082);
nand g499(G1095, G1093, G1094);
nand g500(G1188, G1798, G1805);
not g501(G1900, G1894);
nand g502(G1344, G1894, xenc250);
not g503(G1908, G1902);
nand g504(G1356, G1902, xenc36);
not g505(G1142, G1134);
nand g506(G378, G1234, G1243);
nand g507(G399, G1327, G1330);
not g508(G1331, G1327);
nand g509(G1005, xenc141, G1004);
nand g510(G1015, xenc247, G1014);
not g511(G1764, G1758);
nand g512(G1126, G1758, G1765);
not g513(G1130, G1122);
not g514(G1772, G1766);
nand g515(G1138, G1766, xenc241);
nand g516(G1189, G1187, G1188);
nand g517(G1343, xenc227, xenc181);
nand g518(G1355, G1905, G1908);
nand g519(G324, xenc193, G1098);
not g520(G1099, xenc193);
nand g521(G379, G377, G378);
nand g522(G400, G1322, G1331);
nand g523(G449, G393, G918);
not g524(G1087, xenc105);
nand g525(G1088, xenc105, G1086);
nand g526(G1125, G1761, G1764);
nand g527(G1137, xenc202, G1772);
nand g528(G1345, G1343, G1344);
nand g529(G1357, G1355, G1356);
assign G1397 = G393;
nand g531(G277, G1015, xenc251);
not g532(G1019, G1015);
nand g533(G280, G1005, G1008);
not g534(G1009, G1005);
nand g535(G325, xenc97, G1099);
nand g536(G364, xenc92, G1192);
not g537(G1193, xenc92);
nand g538(G401, G399, G400);
nand g539(G1089, G1078, G1087);
nand g540(G1127, xenc69, G1126);
nand g541(G1139, G1137, G1138);
nand g542(G278, G1010, G1019);
nand g543(G281, G1000, G1009);
nand g544(G326, xenc114, G325);
nand g545(G365, G1184, G1193);
nand g546(G413, G1357, G1360);
not g547(G1361, G1357);
not g548(G1401, xenc32);
nand g549(G445, xenc131, G918);
not g550(G1349, G1345);
nand g551(G1350, G1345, G1348);
assign G1389 = xenc131;
assign G1493 = G449;
assign G1501 = G449;
nand g555(G1689, G1088, xenc100);
nand g556(G279, G277, G278);
nand g557(G282, G280, G281);
nand g558(G346, G1139, xenc151);
not g559(G1143, G1139);
nand g560(G366, G364, xenc2);
nand g561(G414, xenc178, xenc59);
nand g562(G453, G401, G918);
not g563(G1131, G1127);
nand g564(G1132, G1127, G1130);
nand g565(G1351, G1340, G1349);
not g566(G1365, G326);
assign G1405 = G401;
not g568(G285, G279);
nand g569(G347, G1134, G1143);
not g570(G367, xenc89);
nand g571(G415, G413, G414);
not g572(G1393, xenc145);
nand g573(G556, G1501, G1504);
not g574(G1505, G1501);
nand g575(G559, G1493, xenc217);
not g576(G1497, G1493);
not g577(G1693, G1689);
nand g578(G1133, G1122, G1131);
assign G1477 = G445;
assign G1485 = G445;
nand g581(G1809, G1350, G1351);
nand g582(G348, G346, G347);
not g583(G1369, G1365);
not g584(G1409, G1405);
nand g585(G557, G1498, G1505);
nand g586(G560, xenc157, G1497);
assign G1362 = xenc220;
not g588(G1378, G415);
assign G1429 = xenc140;
assign G1437 = xenc140;
assign G1686 = xenc220;
nand g592(G1774, G1132, G1133);
and g593(G1910, xenc55, G853);
and g594(G1918, G856, G367);
nand g595(G544, G1485, G1488);
not g596(G1489, G1485);
nand g597(G547, G1477, xenc126);
not g598(G1481, G1477);
nand g599(G558, G556, G557);
nand g600(G561, G559, G560);
not g601(G1813, G1809);
not g602(G1370, G348);
not g603(G1368, G1362);
nand g604(G417, G1362, G1369);
not g605(G1384, G1378);
nand g606(G424, G1378, G1385);
nand g607(G508, xenc175, xenc252);
not g608(G1441, xenc175);
nand g609(G511, G1429, G1432);
not g610(G1433, G1429);
nand g611(G545, G1482, G1489);
nand g612(G548, G1474, xenc167);
not g613(G564, G558);
not g614(G1692, G1686);
nand g615(G1024, G1686, G1693);
not g616(G1780, G1774);
nand g617(G1148, G1774, xenc50);
not g618(G1916, xenc254);
not g619(G1924, G1918);
nand g620(G416, G1365, G1368);
not g621(G1376, G1370);
nand g622(G421, G1370, G1377);
nand g623(G423, G1381, xenc168);
nand g624(G509, G1434, G1441);
nand g625(G512, xenc64, G1433);
nand g626(G546, G544, G545);
nand g627(G549, G547, G548);
not g628(G719, G561);
assign G722 = G561;
nand g630(G1023, G1689, xenc226);
nand g631(G1147, G1777, G1780);
nand g632(G418, G416, xenc34);
nand g633(G420, xenc7, G1376);
nand g634(G425, G423, G424);
nand g635(G510, G508, G509);
nand g636(G513, xenc215, xenc106);
not g637(G552, G546);
nand g638(G1025, G1023, xenc232);
nand g639(G1149, G1147, G1148);
not g640(G419, xenc113);
nand g641(G422, xenc102, xenc192);
nand g642(G441, G425, G918);
not g643(G516, xenc173);
not g644(G725, xenc117);
assign G728 = xenc117;
not g646(G1029, G1025);
not g647(G1153, G1149);
nand g648(G433, G419, G918);
nand g649(G437, G422, G918);
not g650(G663, xenc104);
assign G666 = xenc104;
and g652(G731, xenc122, G725);
and g653(G746, G722, G725);
and g654(G756, xenc122, G728);
and g655(G770, G722, G728);
assign G1461 = xenc234;
assign G1469 = xenc234;
assign G1413 = G433;
assign G1421 = G433;
assign G1445 = G437;
assign G1453 = G437;
nand g662(G532, G1469, G1472);
not g663(G1473, G1469);
nand g664(G535, G1461, G1464);
not g665(G1465, G1461);
nand g666(G495, G1421, G1424);
not g667(G1425, G1421);
nand g668(G498, G1413, G1416);
not g669(G1417, G1413);
nand g670(G520, G1453, G1456);
not g671(G1457, G1453);
nand g672(G523, xenc162, G1448);
not g673(G1449, xenc162);
nand g674(G533, G1466, G1473);
nand g675(G536, xenc111, G1465);
nand g676(G496, G1418, G1425);
nand g677(G499, G1410, G1417);
nand g678(G521, xenc203, xenc83);
nand g679(G524, xenc121, xenc154);
nand g680(G534, G532, xenc184);
nand g681(G537, G535, xenc187);
nand g682(G497, xenc4, G496);
nand g683(G500, xenc54, G499);
nand g684(G522, G520, G521);
nand g685(G525, G523, G524);
not g686(G540, G534);
not g687(G503, xenc125);
not g688(G528, xenc218);
not g689(G669, G537);
assign G672 = G537;
not g691(G569, G500);
and g692(G588, G566, G500);
not g693(G618, G525);
and g694(G639, G615, G525);
nand g695(G867, xenc231, xenc79, xenc48, G540, G482, xenc244, G503, G487);
assign G588a = G588;
assign G588b = G588;
assign G639a = G639;
assign G639b = G639;
and g700(G675, G663, G669);
and g701(G688, xenc158, G669);
and g702(G696, G663, G672);
and g703(G710, xenc158, G672);
and g704(G73, G949, G867, G932, G932);
and g705(G572, G565, G569);
and g706(G573, G566, G569);
and g707(G621, G614, G618);
and g708(G622, G615, G618);
nand g709(G776, G588a, xenc206, G696, G731, G958);
nand g710(G780, G588a, xenc206, xenc196, xenc27, G958);
nand g711(G784, G588a, xenc206, xenc196, G746, G958);
nand g712(G788, G588a, xenc206, G688, G731, G958);
nand g713(G812, G588b, xenc206, G710, G746, xenc13);
nand g714(G832, G588b, G639b, G696, G770, xenc13);
nand g715(G836, G588b, G639b, G710, xenc27, xenc13);
and g716(G1509, G588a, xenc206, G696, G731, G958);
and g717(G1517, G588a, xenc206, xenc196, xenc27, G958);
and g718(G1525, G588a, xenc206, xenc196, G746, G958);
and g719(G1533, G588a, xenc206, G688, G731, G958);
and g720(G1581, G588b, xenc206, G710, G746, xenc13);
and g721(G1621, G588b, G639b, G696, G770, xenc13);
and g722(G1629, G588b, G639b, G710, xenc27, xenc13);
nand g723(G792, G588a, G622, G696, xenc27, G958);
nand g724(G796, G588b, G622, G696, G746, G958);
nand g725(G800, G588b, G622, G710, G731, G958);
nand g726(G804, G588b, G622, xenc196, G770, G958);
nand g727(G808, G588b, G622, G688, xenc27, xenc13);
nand g728(G816, G573, G639b, G696, xenc27, xenc13);
nand g729(G820, G573, G639b, G696, G746, xenc13);
nand g730(G824, G573, G639b, G710, G731, xenc13);
nand g731(G828, G573, G639b, G688, xenc27, xenc13);
nand g732(G871, G588b, G622, xenc196, G731, xenc245);
nand g733(G873, G573, G639b, xenc196, G731, xenc245);
nand g734(G875, G573, G622, G696, G731, xenc245);
nand g735(G877, G573, G622, xenc196, xenc27, xenc245);
nand g736(G879, G573, G622, xenc196, G746, xenc245);
nand g737(G881, G573, G622, G688, G731, xenc245);
nand g738(G883, G573, G621, xenc196, G731, xenc245);
nand g739(G885, G572, G622, xenc196, G731, xenc245);
and g740(G1541, G588a, G622, G696, xenc27, G958);
and g741(G1549, G588b, G622, G696, G746, G958);
and g742(G1557, G588b, G622, G710, G731, G958);
and g743(G1565, G588b, G622, xenc196, G770, G958);
and g744(G1573, G588b, G622, G688, xenc27, xenc13);
and g745(G1589, G573, G639b, G696, xenc27, xenc13);
and g746(G1597, G573, G639b, G696, G746, xenc13);
and g747(G1605, G573, G639b, G710, G731, xenc13);
and g748(G1613, G573, G639b, G688, xenc27, xenc13);
nand g749(G1, G1509, G1512);
not g750(G1513, G1509);
nand g751(G4, G1517, G1520);
not g752(G1521, G1517);
nand g753(G7, xenc138, G1528);
not g754(G1529, xenc138);
nand g755(G10, G1533, G1536);
not g756(G1537, G1533);
nand g757(G28, G1581, G1584);
not g758(G1585, G1581);
nand g759(G43, G1621, G1624);
not g760(G1625, G1621);
nand g761(G46, G1629, G1632);
not g762(G1633, G1629);
and g763(G886, G871, G873, xenc142, G877, G879, G881, xenc109, G885);
nand g764(G2, G1506, G1513);
nand g765(G5, xenc222, G1521);
nand g766(G8, G1522, G1529);
nand g767(G11, G1530, xenc194);
nand g768(G13, xenc16, G1544);
not g769(G1545, xenc16);
nand g770(G16, xenc94, G1552);
not g771(G1553, xenc94);
nand g772(G19, G1557, xenc165);
not g773(G1561, G1557);
nand g774(G22, G1565, G1568);
not g775(G1569, G1565);
nand g776(G25, G1573, G1576);
not g777(G1577, G1573);
nand g778(G29, xenc63, G1585);
nand g779(G31, G1589, xenc1);
not g780(G1593, G1589);
nand g781(G34, G1597, G1600);
not g782(G1601, G1597);
nand g783(G37, G1605, G1608);
not g784(G1609, G1605);
nand g785(G40, G1613, xenc30);
not g786(G1617, G1613);
nand g787(G44, G1618, G1625);
nand g788(G47, G1626, G1633);
nand g789(G857, xenc135, G780, G784, xenc177, G792, G796, xenc29, xenc164);
nand g790(G860, G808, xenc17, G816, G820, xenc73, xenc45, G832, G836);
and g791(G863, xenc135, G780, G784, xenc177, G792, G796, xenc29, xenc164);
and g792(G865, G808, xenc17, G816, G820, xenc73, xenc45, G832, G836);
nand g793(xenc112, G1, G2);
nand g794(xenc77, G4, G5);
nand g795(G9, G7, G8);
nand g796(G12, G10, G11);
nand g797(G14, xenc87, xenc170);
nand g798(G17, G1546, xenc120);
nand g799(G20, xenc139, G1561);
nand g800(G23, G1562, G1569);
nand g801(G26, G1570, G1577);
nand g802(G30, G28, G29);
nand g803(G32, xenc47, G1593);
nand g804(G35, G1594, G1601);
nand g805(G38, G1602, G1609);
nand g806(G41, G1610, G1617);
nand g807(G45, G43, G44);
nand g808(G48, xenc198, G47);
and g809(G1913, xenc211, G859);
and g810(G1921, G860, G862);
nand g811(G15, xenc153, G14);
nand g812(G18, G16, G17);
nand g813(G21, G19, G20);
nand g814(xenc174, G22, G23);
nand g815(G27, G25, xenc224);
nand g816(G33, G31, G32);
nand g817(G36, G34, G35);
nand g818(xenc49, G37, xenc183);
nand g819(xenc68, G40, G41);
and g820(G887, G863, G865, G886);
nand g821(G462, G863, G865);
and g822(G74, G949, G867, G952, G887);
nand g823(G1637, G1913, G1916);
not g824(G1917, G1913);
nand g825(G1647, G1921, G1924);
not g826(G1925, G1921);
nor g827(G75, xenc201, xenc221);
and g828(G1020, xenc84, G911, G462);
and g829(G1144, G469, G911, G462);
and g830(G1386, G475, G911, G462);
and g831(G1394, G478, G911, G462);
and g832(G1402, G459, G911, G462);
nand g833(G1638, xenc254, G1917);
nand g834(G1648, G1918, G1925);
and g835(G1806, G472, G911, G462);
nand g836(G1639, xenc148, G1638);
nand g837(G1649, G1647, xenc53);
nand g838(G287, G1020, xenc116);
nand g839(G350, G1144, xenc65);
nand g840(G427, G1386, G1393);
nand g841(G429, xenc38, G1401);
nand g842(G431, G1402, G1409);
not g843(G1028, G1020);
not g844(G1152, G1144);
not g845(G1392, G1386);
not g846(G1400, xenc38);
not g847(G1408, G1402);
not g848(G1812, xenc204);
nand g849(G1216, xenc204, G1813);
nand g850(G286, G1025, G1028);
nand g851(G349, G1149, G1152);
nand g852(G426, xenc145, G1392);
nand g853(G428, xenc32, G1400);
nand g854(G430, G1405, G1408);
nand g855(G67, G1639, xenc163);
not g856(G1643, G1639);
nand g857(G70, xenc197, G1652);
not g858(G1653, xenc197);
nand g859(G1215, G1809, G1812);
nand g860(G49, G286, G287);
nand g861(G53, G349, G350);
nand g862(G59, G426, xenc219);
nand g863(G61, G428, G429);
nand g864(G65, G430, G431);
nand g865(G68, G1634, G1643);
nand g866(G71, G1644, G1653);
nand g867(G1217, xenc179, xenc176);
and g868(G51, G49, G50);
and g869(G54, G52, G53);
and g870(xenc152, xenc130, G59);
and g871(G63, G61, G62);
and g872(xenc171, xenc255, xenc242);
nand g873(G69, G67, G68);
nand g874(G72, xenc76, G71);
nand g875(G375, xenc74, xenc150);
not g876(G1221, xenc74);
nand g877(G376, xenc182, G1221);
nand g878(G55, G375, xenc137);
and g879(xenc235, G55, G56);
or g880(xenc0, G1226, keyinput0);
or g881(xenc1, G1592, keyinput1);
and g882(xenc2, G365, keyinput2);
or g883(xenc3, G1211, keyinput3);
or g884(xenc4, G495, keyinput4);
or g885(xenc5, G1822, keyinput5);
and g886(xenc6, G198, keyinput6);
or g887(xenc7, G1373, keyinput7);
or g888(xenc8, G1237, keyinput8);
and g889(xenc9, G1869, keyinput9);
or g890(xenc10, G954, keyinput10);
and g891(xenc11, G1844, keyinput11);
and g892(xenc12, G1732, keyinput12);
and g893(xenc13, G969, keyinput13);
or g894(xenc14, G999, keyinput14);
and g895(xenc15, G1162, keyinput15);
or g896(xenc16, G1541, keyinput16);
and g897(xenc17, G812, keyinput17);
or g898(xenc18, G1673, keyinput18);
or g899(xenc19, G272, keyinput19);
or g900(xenc20, G297, keyinput20);
and g901(xenc21, G1294, keyinput21);
and g902(xenc22, G1662, keyinput22);
or g903(xenc23, G1797, keyinput23);
or g904(xenc24, G1893, keyinput24);
or g905(xenc25, G1260, keyinput25);
or g906(xenc26, G1854, keyinput26);
or g907(xenc27, G756, keyinput27);
and g908(xenc28, G1741, keyinput28);
and g909(xenc29, G800, keyinput29);
or g910(xenc30, G1616, keyinput30);
and g911(xenc31, G1892, keyinput31);
or g912(xenc32, G1397, keyinput32);
or g913(xenc33, G1700, keyinput33);
or g914(xenc34, G417, keyinput34);
and g915(xenc35, G352, keyinput35);
or g916(xenc36, G1909, keyinput36);
or g917(xenc37, G261, keyinput37);
or g918(xenc38, G1394, keyinput38);
and g919(xenc39, G1043, keyinput39);
or g920(xenc40, G956, keyinput40);
or g921(xenc41, G340, keyinput41);
and g922(xenc42, G1326, keyinput42);
or g923(xenc43, G1796, keyinput43);
or g924(xenc44, G1259, keyinput44);
and g925(xenc45, G828, keyinput45);
and g926(xenc46, G1885, keyinput46);
or g927(xenc47, G1586, keyinput47);
and g928(xenc48, G552, keyinput48);
or g929(G39, xenc49, keyinput49);
and g930(xenc50, G1781, keyinput50);
and g931(xenc51, G407, keyinput51);
or g932(xenc52, G1841, keyinput52);
and g933(xenc53, G1648, keyinput53);
or g934(xenc54, G498, keyinput54);
and g935(xenc55, G285, keyinput55);
and g936(xenc56, G404, keyinput56);
and g937(xenc57, G1685, keyinput57);
or g938(xenc58, G1718, keyinput58);
and g939(xenc59, G1361, keyinput59);
and g940(xenc60, G1729, keyinput60);
and g941(xenc61, G302, keyinput61);
and g942(xenc62, G1071, keyinput62);
or g943(xenc63, G1578, keyinput63);
and g944(xenc64, G1426, keyinput64);
or g945(xenc65, G1153, keyinput65);
or g946(xenc66, G1793, keyinput66);
or g947(xenc67, G1061, keyinput67);
and g948(G42, xenc68, keyinput68);
or g949(xenc69, G1125, keyinput69);
or g950(xenc70, G943, keyinput70);
or g951(xenc71, G934, keyinput71);
and g952(xenc72, G202, keyinput72);
or g953(xenc73, G824, keyinput73);
or g954(xenc74, G1217, keyinput74);
or g955(xenc75, G1676, keyinput75);
or g956(xenc76, G70, keyinput76);
or g957(G6, xenc77, keyinput77);
and g958(xenc78, G359, keyinput78);
and g959(xenc79, G564, keyinput79);
and g960(xenc80, G397, keyinput80);
or g961(xenc81, G245, keyinput81);
and g962(xenc82, G296, keyinput82);
or g963(xenc83, G1457, keyinput83);
or g964(xenc84, G457, keyinput84);
or g965(xenc85, G1697, keyinput85);
or g966(xenc86, G1170, keyinput86);
or g967(xenc87, G1538, keyinput87);
or g968(xenc88, G1283, keyinput88);
and g969(xenc89, G366, keyinput89);
and g970(xenc90, G1273, keyinput90);
and g971(xenc91, G1669, keyinput91);
or g972(xenc92, G1189, keyinput92);
and g973(xenc93, G1782, keyinput93);
or g974(xenc94, G1549, keyinput94);
or g975(xenc95, G1750, keyinput95);
and g976(xenc96, G990, keyinput96);
or g977(xenc97, G1090, keyinput97);
and g978(xenc98, G1222, keyinput98);
and g979(xenc99, G1828, keyinput99);
and g980(xenc100, G1089, keyinput100);
or g981(xenc101, G553, keyinput101);
and g982(xenc102, G420, keyinput102);
and g983(xenc103, G358, keyinput103);
and g984(xenc104, G513, keyinput104);
or g985(xenc105, G1083, keyinput105);
or g986(xenc106, G512, keyinput106);
and g987(xenc107, G1312, keyinput107);
and g988(xenc108, G1726, keyinput108);
and g989(xenc109, G883, keyinput109);
and g990(xenc110, G305, keyinput110);
and g991(xenc111, G1458, keyinput111);
or g992(G3, xenc112, keyinput112);
and g993(xenc113, G418, keyinput113);
or g994(xenc114, G324, keyinput114);
and g995(xenc115, G1785, keyinput115);
or g996(xenc116, G1029, keyinput116);
and g997(xenc117, G549, keyinput117);
and g998(xenc118, G1335, keyinput118);
and g999(xenc119, G1174, keyinput119);
and g1000(xenc120, G1553, keyinput120);
and g1001(xenc121, G1442, keyinput121);
and g1002(xenc122, G719, keyinput122);
or g1003(xenc123, G1309, keyinput123);
and g1004(xenc124, G1724, keyinput124);
and g1005(xenc125, G497, keyinput125);
and g1006(xenc126, G1480, keyinput126);
and g1007(xenc127, G1860, keyinput127);
or g1008(xenc128, G318, keyinput128);
and g1009(xenc129, G1171, keyinput129);
or g1010(xenc130, G58, keyinput130);
or g1011(xenc131, G379, keyinput131);
or g1012(xenc132, G1804, keyinput132);
or g1013(xenc133, G1325, keyinput133);
or g1014(xenc134, G1166, keyinput134);
and g1015(xenc135, G776, keyinput135);
and g1016(xenc136, G385, keyinput136);
and g1017(xenc137, G376, keyinput137);
and g1018(xenc138, G1525, keyinput138);
and g1019(xenc139, G1554, keyinput139);
and g1020(xenc140, G453, keyinput140);
and g1021(xenc141, G1003, keyinput141);
and g1022(xenc142, G875, keyinput142);
or g1023(xenc143, G1165, keyinput143);
and g1024(xenc144, G1183, keyinput144);
or g1025(xenc145, G1389, keyinput145);
and g1026(xenc146, G1038, keyinput146);
or g1027(xenc147, G179, keyinput147);
or g1028(xenc148, G1637, keyinput148);
and g1029(xenc149, G1657, keyinput149);
or g1030(xenc150, G1220, keyinput150);
or g1031(xenc151, G1142, keyinput151);
and g1032(G60, xenc152, keyinput152);
and g1033(xenc153, G13, keyinput153);
or g1034(xenc154, G1449, keyinput154);
and g1035(xenc155, G310, keyinput155);
and g1036(xenc156, G1249, keyinput156);
or g1037(xenc157, G1490, keyinput157);
or g1038(xenc158, G666, keyinput158);
or g1039(xenc159, G1833, keyinput159);
and g1040(xenc160, G1338, keyinput160);
and g1041(xenc161, G262, keyinput161);
and g1042(xenc162, G1445, keyinput162);
or g1043(xenc163, G1642, keyinput163);
or g1044(xenc164, G804, keyinput164);
or g1045(xenc165, G1560, keyinput165);
or g1046(xenc166, G1117, keyinput166);
or g1047(xenc167, G1481, keyinput167);
or g1048(xenc168, G1384, keyinput168);
or g1049(xenc169, G355, keyinput169);
or g1050(xenc170, G1545, keyinput170);
and g1051(G66, xenc171, keyinput171);
or g1052(xenc172, G1121, keyinput172);
or g1053(xenc173, G510, keyinput173);
or g1054(G24, xenc174, keyinput174);
or g1055(xenc175, G1437, keyinput175);
and g1056(xenc176, G1216, keyinput176);
or g1057(xenc177, G788, keyinput177);
and g1058(xenc178, G1352, keyinput178);
or g1059(xenc179, G1215, keyinput179);
or g1060(xenc180, G1303, keyinput180);
and g1061(xenc181, G1900, keyinput181);
and g1062(xenc182, G1212, keyinput182);
or g1063(xenc183, G38, keyinput183);
and g1064(xenc184, G533, keyinput184);
or g1065(xenc185, G335, keyinput185);
and g1066(xenc186, G492, keyinput186);
and g1067(xenc187, G536, keyinput187);
or g1068(xenc188, G360, keyinput188);
or g1069(xenc189, G1244, keyinput189);
or g1070(xenc190, G1239, keyinput190);
or g1071(xenc191, G257, keyinput191);
or g1072(xenc192, G421, keyinput192);
or g1073(xenc193, G1095, keyinput193);
and g1074(xenc194, G1537, keyinput194);
and g1075(xenc195, G1281, keyinput195);
and g1076(xenc196, G675, keyinput196);
and g1077(xenc197, G1649, keyinput197);
or g1078(xenc198, G46, keyinput198);
or g1079(xenc199, G1316, keyinput199);
or g1080(xenc200, G1740, keyinput200);
and g1081(xenc201, G73, keyinput201);
or g1082(xenc202, G1769, keyinput202);
or g1083(xenc203, G1450, keyinput203);
or g1084(xenc204, G1806, keyinput204);
or g1085(xenc205, G1717, keyinput205);
and g1086(xenc206, G639a, keyinput206);
or g1087(xenc207, G388, keyinput207);
and g1088(xenc208, G1665, keyinput208);
or g1089(xenc209, G398, keyinput209);
and g1090(xenc210, G1708, keyinput210);
and g1091(xenc211, G857, keyinput211);
or g1092(xenc212, G241, keyinput212);
and g1093(xenc213, G274, keyinput213);
or g1094(xenc214, G1339, keyinput214);
or g1095(xenc215, G511, keyinput215);
and g1096(xenc216, G1164, keyinput216);
or g1097(xenc217, G1496, keyinput217);
or g1098(xenc218, G522, keyinput218);
or g1099(xenc219, G427, keyinput219);
and g1100(xenc220, G282, keyinput220);
and g1101(xenc221, G74, keyinput221);
and g1102(xenc222, G1514, keyinput222);
or g1103(xenc223, G907, keyinput223);
or g1104(xenc224, G26, keyinput224);
and g1105(xenc225, G1050, keyinput225);
or g1106(xenc226, G1692, keyinput226);
or g1107(xenc227, G1897, keyinput227);
and g1108(xenc228, G1230, keyinput228);
and g1109(xenc229, G1110, keyinput229);
and g1110(xenc230, G1721, keyinput230);
and g1111(xenc231, G516, keyinput231);
and g1112(xenc232, G1024, keyinput232);
and g1113(xenc233, G988, keyinput233);
or g1114(xenc234, G441, keyinput234);
or g1115(G57, xenc235, keyinput235);
or g1116(xenc236, G1862, keyinput236);
or g1117(xenc237, G1830, keyinput237);
and g1118(xenc238, G1289, keyinput238);
or g1119(xenc239, G1207, keyinput239);
and g1120(xenc240, G1677, keyinput240);
and g1121(xenc241, G1773, keyinput241);
or g1122(xenc242, G65, keyinput242);
or g1123(xenc243, G1876, keyinput243);
or g1124(xenc244, G528, keyinput244);
or g1125(xenc245, G979, keyinput245);
and g1126(xenc246, G1293, keyinput246);
or g1127(xenc247, G1013, keyinput247);
and g1128(xenc248, G1710, keyinput248);
or g1129(xenc249, G390, keyinput249);
and g1130(xenc250, G1901, keyinput250);
or g1131(xenc251, G1018, keyinput251);
or g1132(xenc252, G1440, keyinput252);
and g1133(xenc253, G392, keyinput253);
and g1134(xenc254, G1910, keyinput254);
and g1135(xenc255, G64, keyinput255);
endmodule
