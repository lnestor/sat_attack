
module c3540 ( N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, 
        N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, 
        N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, 
        N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, 
        N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, 
        N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, 
        N5231, N5360, N5361, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31 );
  input N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116,
         N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190,
         N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264,
         N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330,
         N343, N349, N350, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31;
  output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815,
         N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231,
         N5360, N5361;
  wire   n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971;

  MUX21X1 U494 ( .IN1(n480), .IN2(n481), .S(n482), .Q(N5361) );
  XNOR2X1 U495 ( .IN1(n483), .IN2(n484), .Q(n482) );
  AOI21X1 U496 ( .IN1(N5120), .IN2(N5102), .IN3(n485), .QN(n484) );
  NAND2X0 U497 ( .IN1(n480), .IN2(keyinput31), .QN(n481) );
  XNOR2X1 U498 ( .IN1(n486), .IN2(keyinput30), .Q(n480) );
  XOR2X1 U499 ( .IN1(n487), .IN2(n486), .Q(N5360) );
  XOR3X1 U500 ( .IN1(N4815), .IN2(N5045), .IN3(n488), .Q(n486) );
  XNOR2X1 U501 ( .IN1(N5078), .IN2(N5047), .Q(n488) );
  MUX21X1 U502 ( .IN1(n483), .IN2(n489), .S(n490), .Q(n487) );
  XOR2X1 U503 ( .IN1(n491), .IN2(n492), .Q(n490) );
  MUX21X1 U504 ( .IN1(N5120), .IN2(N350), .S(n493), .Q(n492) );
  NOR2X0 U505 ( .IN1(n493), .IN2(n494), .QN(n491) );
  INVX0 U506 ( .INP(N5102), .ZN(n494) );
  AND2X1 U507 ( .IN1(N213), .IN2(n495), .Q(n493) );
  NOR2X0 U508 ( .IN1(n496), .IN2(n497), .QN(n489) );
  INVX0 U509 ( .INP(n498), .ZN(n497) );
  NAND2X0 U510 ( .IN1(n499), .IN2(n498), .QN(n483) );
  NAND2X0 U511 ( .IN1(n500), .IN2(N5121), .QN(n498) );
  XOR2X1 U512 ( .IN1(keyinput29), .IN2(n496), .Q(n499) );
  NOR2X0 U513 ( .IN1(n500), .IN2(N5121), .QN(n496) );
  NAND3X0 U514 ( .IN1(n501), .IN2(N5192), .IN3(N213), .QN(N5231) );
  NAND2X0 U515 ( .IN1(n485), .IN2(n495), .QN(n501) );
  NAND4X0 U516 ( .IN1(n502), .IN2(n500), .IN3(n485), .IN4(n503), .QN(N5192) );
  NOR4X0 U517 ( .IN1(N5121), .IN2(N5078), .IN3(N5047), .IN4(N5045), .QN(n503)
         );
  NOR2X0 U518 ( .IN1(N5102), .IN2(N5120), .QN(n485) );
  AO222X1 U519 ( .IN1(n504), .IN2(n505), .IN3(n506), .IN4(n507), .IN5(n508), 
        .IN6(n509), .Q(N5121) );
  AOI222X1 U520 ( .IN1(n510), .IN2(n511), .IN3(n512), .IN4(n513), .IN5(n514), 
        .IN6(n515), .QN(n507) );
  OA221X1 U521 ( .IN1(n516), .IN2(n517), .IN3(n518), .IN4(n519), .IN5(n520), 
        .Q(n515) );
  OA222X1 U522 ( .IN1(n521), .IN2(n522), .IN3(n523), .IN4(n524), .IN5(n525), 
        .IN6(n526), .Q(n520) );
  XNOR2X1 U523 ( .IN1(keyinput13), .IN2(n527), .Q(n524) );
  OA221X1 U524 ( .IN1(n528), .IN2(n529), .IN3(n530), .IN4(n531), .IN5(n532), 
        .Q(n514) );
  OA21X1 U525 ( .IN1(n533), .IN2(n534), .IN3(n535), .Q(n532) );
  OA221X1 U526 ( .IN1(n530), .IN2(n536), .IN3(n516), .IN4(n537), .IN5(n538), 
        .Q(n511) );
  OA222X1 U527 ( .IN1(n518), .IN2(n539), .IN3(n525), .IN4(n540), .IN5(n521), 
        .IN6(n541), .Q(n538) );
  OA221X1 U528 ( .IN1(n527), .IN2(n542), .IN3(n528), .IN4(n543), .IN5(n544), 
        .Q(n510) );
  OA21X1 U529 ( .IN1(n533), .IN2(n545), .IN3(n546), .Q(n544) );
  OA21X1 U530 ( .IN1(n547), .IN2(n548), .IN3(n549), .Q(n506) );
  XNOR2X1 U531 ( .IN1(n550), .IN2(n551), .Q(n504) );
  AND2X1 U532 ( .IN1(n552), .IN2(n553), .Q(n551) );
  AO21X1 U533 ( .IN1(n554), .IN2(n555), .IN3(n556), .Q(N5120) );
  OA221X1 U534 ( .IN1(N50), .IN2(n557), .IN3(n558), .IN4(n559), .IN5(n560), 
        .Q(n556) );
  OA21X1 U535 ( .IN1(n548), .IN2(n561), .IN3(n549), .Q(n560) );
  MUX21X1 U536 ( .IN1(N50), .IN2(n562), .S(n563), .Q(n559) );
  MUX21X1 U537 ( .IN1(n564), .IN2(n565), .S(n566), .Q(n562) );
  NAND4X0 U538 ( .IN1(n567), .IN2(n568), .IN3(n569), .IN4(n570), .QN(n565) );
  OA221X1 U539 ( .IN1(n530), .IN2(n542), .IN3(n516), .IN4(n545), .IN5(n571), 
        .Q(n570) );
  OA22X1 U540 ( .IN1(n525), .IN2(n572), .IN3(n518), .IN4(n540), .Q(n571) );
  AOI22X1 U541 ( .IN1(N124), .IN2(n573), .IN3(N143), .IN4(n574), .QN(n569) );
  NAND2X0 U542 ( .IN1(N137), .IN2(n575), .QN(n568) );
  XOR2X1 U543 ( .IN1(n576), .IN2(keyinput16), .Q(n567) );
  NAND2X0 U544 ( .IN1(N128), .IN2(n577), .QN(n576) );
  NAND4X0 U545 ( .IN1(n578), .IN2(n579), .IN3(n580), .IN4(n581), .QN(n564) );
  OA22X1 U546 ( .IN1(n582), .IN2(n519), .IN3(n521), .IN4(n534), .Q(n581) );
  XNOR2X1 U547 ( .IN1(n583), .IN2(keyinput12), .Q(n582) );
  OA22X1 U548 ( .IN1(n523), .IN2(n518), .IN3(n516), .IN4(n513), .Q(n580) );
  OA22X1 U549 ( .IN1(n530), .IN2(n536), .IN3(n522), .IN4(n528), .Q(n579) );
  OA22X1 U550 ( .IN1(n527), .IN2(n531), .IN3(n517), .IN4(n533), .Q(n578) );
  AO21X1 U551 ( .IN1(n505), .IN2(n584), .IN3(n509), .Q(n555) );
  AO21X1 U552 ( .IN1(n585), .IN2(n508), .IN3(n586), .Q(n584) );
  XNOR2X1 U553 ( .IN1(n561), .IN2(n587), .Q(n554) );
  NOR2X0 U554 ( .IN1(n588), .IN2(n589), .QN(n587) );
  INVX0 U555 ( .INP(n590), .ZN(n588) );
  XOR2X1 U556 ( .IN1(n591), .IN2(n592), .Q(n561) );
  NAND2X0 U557 ( .IN1(n593), .IN2(n594), .QN(n591) );
  INVX0 U558 ( .INP(n595), .ZN(n593) );
  NAND2X0 U559 ( .IN1(n596), .IN2(n597), .QN(N5078) );
  NAND3X0 U560 ( .IN1(n549), .IN2(n598), .IN3(n599), .QN(n597) );
  AOI222X1 U561 ( .IN1(n600), .IN2(n601), .IN3(n602), .IN4(n603), .IN5(n604), 
        .IN6(n605), .QN(n599) );
  OA221X1 U562 ( .IN1(n530), .IN2(n534), .IN3(n519), .IN4(n516), .IN5(n606), 
        .Q(n605) );
  OA222X1 U563 ( .IN1(n518), .IN2(n529), .IN3(n525), .IN4(n607), .IN5(n521), 
        .IN6(n608), .Q(n606) );
  OA221X1 U564 ( .IN1(n527), .IN2(n522), .IN3(n528), .IN4(n609), .IN5(n610), 
        .Q(n604) );
  OA21X1 U565 ( .IN1(n526), .IN2(n533), .IN3(n535), .Q(n610) );
  AO221X1 U566 ( .IN1(n611), .IN2(n523), .IN3(n612), .IN4(n613), .IN5(n614), 
        .Q(n603) );
  OA221X1 U567 ( .IN1(n517), .IN2(n530), .IN3(n516), .IN4(n531), .IN5(n615), 
        .Q(n601) );
  OA222X1 U568 ( .IN1(n518), .IN2(n537), .IN3(n525), .IN4(n545), .IN5(n521), 
        .IN6(n542), .Q(n615) );
  OA221X1 U569 ( .IN1(n527), .IN2(n513), .IN3(n528), .IN4(n539), .IN5(n616), 
        .Q(n600) );
  OA21X1 U570 ( .IN1(n533), .IN2(n536), .IN3(n546), .Q(n616) );
  NAND2X0 U571 ( .IN1(n617), .IN2(n618), .QN(n598) );
  MUX21X1 U572 ( .IN1(n619), .IN2(n620), .S(n621), .Q(n596) );
  OA21X1 U573 ( .IN1(n622), .IN2(n623), .IN3(n624), .Q(n620) );
  NAND2X0 U574 ( .IN1(n625), .IN2(n622), .QN(n619) );
  AO221X1 U575 ( .IN1(n626), .IN2(n505), .IN3(n585), .IN4(n509), .IN5(n627), 
        .Q(N5102) );
  NOR3X0 U576 ( .IN1(n628), .IN2(n629), .IN3(n630), .QN(n627) );
  XOR2X1 U577 ( .IN1(n631), .IN2(keyinput24), .Q(n629) );
  OR2X1 U578 ( .IN1(n632), .IN2(n548), .Q(n631) );
  AO222X1 U579 ( .IN1(n633), .IN2(n634), .IN3(n512), .IN4(n536), .IN5(n635), 
        .IN6(n636), .Q(n628) );
  OA221X1 U580 ( .IN1(n530), .IN2(n537), .IN3(n516), .IN4(n542), .IN5(n637), 
        .Q(n636) );
  OA222X1 U581 ( .IN1(n518), .IN2(n541), .IN3(n525), .IN4(n543), .IN5(n521), 
        .IN6(n540), .Q(n637) );
  INVX0 U582 ( .INP(N128), .ZN(n543) );
  OA221X1 U583 ( .IN1(n527), .IN2(n545), .IN3(n528), .IN4(n572), .IN5(n638), 
        .Q(n635) );
  OA21X1 U584 ( .IN1(n533), .IN2(n539), .IN3(n546), .Q(n638) );
  INVX0 U585 ( .INP(N125), .ZN(n572) );
  OA221X1 U586 ( .IN1(n530), .IN2(n513), .IN3(n516), .IN4(n531), .IN5(n639), 
        .Q(n634) );
  OA222X1 U587 ( .IN1(n518), .IN2(n534), .IN3(n525), .IN4(n522), .IN5(n521), 
        .IN6(n519), .Q(n639) );
  OA221X1 U588 ( .IN1(n527), .IN2(n517), .IN3(n526), .IN4(n528), .IN5(n640), 
        .Q(n633) );
  OA21X1 U589 ( .IN1(n523), .IN2(n533), .IN3(n535), .Q(n640) );
  XNOR3X1 U590 ( .IN1(keyinput28), .IN2(n585), .IN3(n641), .Q(n626) );
  NAND2X0 U591 ( .IN1(n550), .IN2(n508), .QN(n641) );
  NAND2X0 U592 ( .IN1(n642), .IN2(n552), .QN(n508) );
  NAND2X0 U593 ( .IN1(n643), .IN2(n644), .QN(n552) );
  XOR2X1 U594 ( .IN1(n553), .IN2(keyinput26), .Q(n642) );
  AO21X1 U595 ( .IN1(n644), .IN2(n645), .IN3(n643), .Q(n553) );
  NAND2X0 U596 ( .IN1(n646), .IN2(n647), .QN(n645) );
  XNOR2X1 U597 ( .IN1(n648), .IN2(keyinput25), .Q(n644) );
  OR2X1 U598 ( .IN1(n647), .IN2(n646), .Q(n648) );
  INVX0 U599 ( .INP(n547), .ZN(n646) );
  INVX0 U600 ( .INP(n586), .ZN(n550) );
  AO21X1 U601 ( .IN1(n649), .IN2(n650), .IN3(n651), .Q(n586) );
  XNOR2X1 U602 ( .IN1(n632), .IN2(n652), .Q(n585) );
  AOI21X1 U603 ( .IN1(n547), .IN2(n643), .IN3(n653), .QN(n652) );
  NAND2X0 U604 ( .IN1(n654), .IN2(n655), .QN(N5047) );
  NAND4X0 U605 ( .IN1(n656), .IN2(n657), .IN3(n658), .IN4(n659), .QN(n655) );
  OA21X1 U606 ( .IN1(n660), .IN2(n661), .IN3(n549), .Q(n659) );
  OA221X1 U607 ( .IN1(N107), .IN2(n662), .IN3(n663), .IN4(n664), .IN5(n665), 
        .Q(n660) );
  NAND3X0 U608 ( .IN1(n666), .IN2(n667), .IN3(n612), .QN(n665) );
  NAND4X0 U609 ( .IN1(n663), .IN2(N58), .IN3(n668), .IN4(n669), .QN(n667) );
  INVX0 U610 ( .INP(n670), .ZN(n669) );
  NOR2X0 U611 ( .IN1(N50), .IN2(N45), .QN(n668) );
  XOR2X1 U612 ( .IN1(keyinput19), .IN2(n671), .Q(n666) );
  NOR2X0 U613 ( .IN1(n672), .IN2(n673), .QN(n671) );
  INVX0 U614 ( .INP(n674), .ZN(n663) );
  NAND4X0 U615 ( .IN1(n535), .IN2(n675), .IN3(n676), .IN4(n677), .QN(n658) );
  OA221X1 U616 ( .IN1(n519), .IN2(n530), .IN3(n522), .IN4(n516), .IN5(n678), 
        .Q(n677) );
  OA222X1 U617 ( .IN1(n518), .IN2(n608), .IN3(n525), .IN4(n609), .IN5(n521), 
        .IN6(n607), .Q(n678) );
  INVX0 U618 ( .INP(N317), .ZN(n607) );
  INVX0 U619 ( .INP(N322), .ZN(n609) );
  AOI22X1 U620 ( .IN1(n573), .IN2(N326), .IN3(n574), .IN4(N294), .QN(n676) );
  NAND2X0 U621 ( .IN1(n575), .IN2(N303), .QN(n675) );
  NAND2X0 U622 ( .IN1(n679), .IN2(n617), .QN(n657) );
  NAND4X0 U623 ( .IN1(n546), .IN2(n680), .IN3(n681), .IN4(n682), .QN(n656) );
  OA221X1 U624 ( .IN1(n523), .IN2(n530), .IN3(n516), .IN4(n517), .IN5(n683), 
        .Q(n682) );
  OA222X1 U625 ( .IN1(n518), .IN2(n536), .IN3(n684), .IN4(n542), .IN5(n521), 
        .IN6(n537), .Q(n683) );
  XNOR2X1 U626 ( .IN1(n583), .IN2(keyinput11), .Q(n684) );
  OA22X1 U627 ( .IN1(n528), .IN2(n545), .IN3(n527), .IN4(n531), .Q(n681) );
  NAND2X0 U628 ( .IN1(N68), .IN2(n575), .QN(n680) );
  INVX0 U629 ( .INP(n533), .ZN(n575) );
  MUX21X1 U630 ( .IN1(n685), .IN2(n624), .S(n622), .Q(n654) );
  OA21X1 U631 ( .IN1(n623), .IN2(n686), .IN3(n687), .Q(n624) );
  INVX0 U632 ( .INP(n625), .ZN(n685) );
  AO222X1 U633 ( .IN1(n688), .IN2(n689), .IN3(n690), .IN4(n691), .IN5(n692), 
        .IN6(n693), .Q(N5045) );
  NAND2X0 U634 ( .IN1(n687), .IN2(n694), .QN(n693) );
  NAND3X0 U635 ( .IN1(n622), .IN2(n625), .IN3(n621), .QN(n694) );
  XOR2X1 U636 ( .IN1(n695), .IN2(n618), .Q(n621) );
  NOR2X0 U637 ( .IN1(n696), .IN2(n623), .QN(n625) );
  XOR2X1 U638 ( .IN1(n697), .IN2(n679), .Q(n622) );
  INVX0 U639 ( .INP(n509), .ZN(n687) );
  XNOR2X1 U640 ( .IN1(keyinput27), .IN2(n689), .Q(n692) );
  OA221X1 U641 ( .IN1(n698), .IN2(n699), .IN3(n700), .IN4(n701), .IN5(n702), 
        .Q(n691) );
  NAND4X0 U642 ( .IN1(n546), .IN2(n703), .IN3(n704), .IN4(n705), .QN(n702) );
  OA221X1 U643 ( .IN1(n528), .IN2(n541), .IN3(n516), .IN4(n513), .IN5(n706), 
        .Q(n705) );
  OA222X1 U644 ( .IN1(n518), .IN2(n542), .IN3(n525), .IN4(n539), .IN5(n521), 
        .IN6(n545), .Q(n706) );
  OA22X1 U645 ( .IN1(n527), .IN2(n536), .IN3(n533), .IN4(n537), .Q(n704) );
  XOR2X1 U646 ( .IN1(keyinput17), .IN2(n707), .Q(n703) );
  NOR2X0 U647 ( .IN1(n530), .IN2(n531), .QN(n707) );
  AO221X1 U648 ( .IN1(N317), .IN2(n573), .IN3(N116), .IN4(n574), .IN5(n708), 
        .Q(n701) );
  OAI21X1 U649 ( .IN1(n533), .IN2(n522), .IN3(n535), .QN(n708) );
  AO221X1 U650 ( .IN1(N107), .IN2(n709), .IN3(n710), .IN4(N97), .IN5(n711), 
        .Q(n700) );
  AO222X1 U651 ( .IN1(N303), .IN2(n577), .IN3(N311), .IN4(n583), .IN5(n712), 
        .IN6(N294), .Q(n711) );
  XNOR2X1 U652 ( .IN1(n602), .IN2(keyinput9), .Q(n699) );
  OA221X1 U653 ( .IN1(n713), .IN2(n714), .IN3(N87), .IN4(n662), .IN5(n664), 
        .Q(n698) );
  OA21X1 U654 ( .IN1(n715), .IN2(n716), .IN3(n549), .Q(n690) );
  XNOR2X1 U655 ( .IN1(n716), .IN2(n717), .Q(n689) );
  OA22X1 U656 ( .IN1(n695), .IN2(n618), .IN3(n718), .IN4(n719), .Q(n717) );
  XOR2X1 U657 ( .IN1(n720), .IN2(n721), .Q(n618) );
  NAND2X0 U658 ( .IN1(n718), .IN2(n722), .QN(n720) );
  XOR2X1 U659 ( .IN1(n723), .IN2(n724), .Q(n716) );
  AND2X1 U660 ( .IN1(n725), .IN2(n718), .Q(n724) );
  NOR2X0 U661 ( .IN1(n686), .IN2(n623), .QN(n688) );
  AO21X1 U662 ( .IN1(n726), .IN2(n727), .IN3(n728), .Q(N5002) );
  MUX21X1 U663 ( .IN1(n729), .IN2(n730), .S(n731), .Q(n728) );
  NOR2X0 U664 ( .IN1(n726), .IN2(n732), .QN(n730) );
  XOR3X1 U665 ( .IN1(n589), .IN2(n651), .IN3(n733), .Q(n732) );
  MUX21X1 U666 ( .IN1(n734), .IN2(n590), .S(n735), .Q(n733) );
  NAND3X0 U667 ( .IN1(n632), .IN2(n547), .IN3(n643), .QN(n590) );
  AND2X1 U668 ( .IN1(n649), .IN2(n736), .Q(n643) );
  NAND2X0 U669 ( .IN1(n649), .IN2(n737), .QN(n734) );
  NAND3X0 U670 ( .IN1(n547), .IN2(n736), .IN3(n632), .QN(n737) );
  AO21X1 U671 ( .IN1(n650), .IN2(n738), .IN3(n739), .Q(n651) );
  AO22X1 U672 ( .IN1(n740), .IN2(n595), .IN3(n632), .IN4(n653), .Q(n589) );
  AO22X1 U673 ( .IN1(n741), .IN2(n742), .IN3(n547), .IN4(n647), .Q(n653) );
  AO21X1 U674 ( .IN1(n743), .IN2(n742), .IN3(n744), .Q(n647) );
  XNOR2X1 U675 ( .IN1(n745), .IN2(n746), .Q(n547) );
  NAND2X0 U676 ( .IN1(n718), .IN2(n747), .QN(n745) );
  XOR2X1 U677 ( .IN1(n748), .IN2(n749), .Q(n632) );
  NOR2X0 U678 ( .IN1(n750), .IN2(n595), .QN(n749) );
  OA21X1 U679 ( .IN1(n751), .IN2(n752), .IN3(N116), .Q(n729) );
  XOR2X1 U680 ( .IN1(n753), .IN2(keyinput3), .Q(n752) );
  NAND2X0 U681 ( .IN1(N97), .IN2(n534), .QN(n753) );
  NOR2X0 U682 ( .IN1(N97), .IN2(n534), .QN(n751) );
  AO21X1 U683 ( .IN1(n670), .IN2(n536), .IN3(n754), .Q(n727) );
  MUX21X1 U684 ( .IN1(n537), .IN2(n755), .S(n513), .Q(n754) );
  NOR2X0 U685 ( .IN1(n531), .IN2(n756), .QN(n755) );
  NOR2X0 U686 ( .IN1(n513), .IN2(n531), .QN(n670) );
  INVX0 U687 ( .INP(n500), .ZN(N4944) );
  MUX21X1 U688 ( .IN1(n757), .IN2(n758), .S(n630), .Q(n500) );
  XNOR2X1 U689 ( .IN1(n649), .IN2(n759), .Q(n758) );
  AOI21X1 U690 ( .IN1(n760), .IN2(n761), .IN3(n744), .QN(n759) );
  NOR2X0 U691 ( .IN1(n760), .IN2(n761), .QN(n744) );
  INVX0 U692 ( .INP(n736), .ZN(n761) );
  AO221X1 U693 ( .IN1(n762), .IN2(n763), .IN3(n764), .IN4(n765), .IN5(n766), 
        .Q(n757) );
  AO22X1 U694 ( .IN1(n767), .IN2(n768), .IN3(n512), .IN4(n531), .Q(n766) );
  INVX0 U695 ( .INP(n557), .ZN(n512) );
  NAND2X0 U696 ( .IN1(n548), .IN2(n558), .QN(n557) );
  OA221X1 U697 ( .IN1(n517), .IN2(n530), .IN3(n523), .IN4(n516), .IN5(n769), 
        .Q(n768) );
  OA222X1 U698 ( .IN1(n522), .IN2(n518), .IN3(n525), .IN4(n529), .IN5(n526), 
        .IN6(n521), .Q(n769) );
  OA221X1 U699 ( .IN1(n527), .IN2(n534), .IN3(n528), .IN4(n608), .IN5(n770), 
        .Q(n767) );
  OA21X1 U700 ( .IN1(n519), .IN2(n533), .IN3(n535), .Q(n770) );
  XNOR2X1 U701 ( .IN1(n736), .IN2(keyinput23), .Q(n764) );
  XNOR2X1 U702 ( .IN1(n771), .IN2(n772), .Q(n736) );
  NAND2X0 U703 ( .IN1(n718), .IN2(n773), .QN(n771) );
  OA221X1 U704 ( .IN1(n530), .IN2(n513), .IN3(n516), .IN4(n536), .IN5(n774), 
        .Q(n763) );
  OA222X1 U705 ( .IN1(n518), .IN2(n545), .IN3(n525), .IN4(n541), .IN5(n521), 
        .IN6(n539), .Q(n774) );
  INVX0 U706 ( .INP(N143), .ZN(n539) );
  INVX0 U707 ( .INP(N137), .ZN(n541) );
  INVX0 U708 ( .INP(N150), .ZN(n545) );
  OA221X1 U709 ( .IN1(n527), .IN2(n537), .IN3(n528), .IN4(n540), .IN5(n775), 
        .Q(n762) );
  OA21X1 U710 ( .IN1(n533), .IN2(n542), .IN3(n546), .Q(n775) );
  INVX0 U711 ( .INP(N132), .ZN(n540) );
  INVX0 U712 ( .INP(n502), .ZN(N4815) );
  MUX21X1 U713 ( .IN1(n776), .IN2(n777), .S(n630), .Q(n502) );
  INVX0 U714 ( .INP(n549), .ZN(n630) );
  NOR2X0 U715 ( .IN1(n509), .IN2(n505), .QN(n549) );
  INVX0 U716 ( .INP(n623), .ZN(n505) );
  NAND2X0 U717 ( .IN1(N1), .IN2(n778), .QN(n509) );
  NAND3X0 U718 ( .IN1(N13), .IN2(n779), .IN3(N45), .QN(n778) );
  XNOR2X1 U719 ( .IN1(N330), .IN2(n780), .Q(n777) );
  NAND4X0 U720 ( .IN1(n781), .IN2(n782), .IN3(n783), .IN4(n784), .QN(n776) );
  NAND4X0 U721 ( .IN1(n535), .IN2(n785), .IN3(n786), .IN4(n787), .QN(n784) );
  AOI221X1 U722 ( .IN1(n710), .IN2(N283), .IN3(N329), .IN4(n573), .IN5(n788), 
        .QN(n787) );
  AO222X1 U723 ( .IN1(N322), .IN2(n577), .IN3(N326), .IN4(n583), .IN5(N317), 
        .IN6(n712), .Q(n788) );
  INVX0 U724 ( .INP(n525), .ZN(n583) );
  INVX0 U725 ( .INP(n521), .ZN(n577) );
  INVX0 U726 ( .INP(n528), .ZN(n573) );
  INVX0 U727 ( .INP(n530), .ZN(n710) );
  OA22X1 U728 ( .IN1(n527), .IN2(n529), .IN3(n533), .IN4(n608), .Q(n786) );
  INVX0 U729 ( .INP(N311), .ZN(n608) );
  INVX0 U730 ( .INP(N303), .ZN(n529) );
  XOR2X1 U731 ( .IN1(keyinput18), .IN2(n789), .Q(n785) );
  NOR2X0 U732 ( .IN1(n790), .IN2(n526), .QN(n789) );
  INVX0 U733 ( .INP(N294), .ZN(n526) );
  XNOR2X1 U734 ( .IN1(n709), .IN2(keyinput14), .Q(n790) );
  INVX0 U735 ( .INP(n516), .ZN(n709) );
  NOR2X0 U736 ( .IN1(n566), .IN2(n558), .QN(n535) );
  NAND2X0 U737 ( .IN1(n602), .IN2(n791), .QN(n783) );
  AO222X1 U738 ( .IN1(n792), .IN2(n519), .IN3(n793), .IN4(n612), .IN5(n614), 
        .IN6(N1947), .Q(n791) );
  MUX21X1 U739 ( .IN1(n794), .IN2(n795), .S(n672), .Q(n793) );
  XNOR2X1 U740 ( .IN1(keyinput6), .IN2(n662), .Q(n792) );
  INVX0 U741 ( .INP(n611), .ZN(n662) );
  NOR2X0 U742 ( .IN1(n614), .IN2(n612), .QN(n611) );
  INVX0 U743 ( .INP(n714), .ZN(n612) );
  NAND2X0 U744 ( .IN1(N33), .IN2(n796), .QN(n714) );
  INVX0 U745 ( .INP(n664), .ZN(n614) );
  NAND2X0 U746 ( .IN1(n796), .IN2(n566), .QN(n664) );
  INVX0 U747 ( .INP(n661), .ZN(n602) );
  NAND2X0 U748 ( .IN1(n715), .IN2(n558), .QN(n661) );
  NAND4X0 U749 ( .IN1(n546), .IN2(n797), .IN3(n798), .IN4(n799), .QN(n782) );
  OA221X1 U750 ( .IN1(n531), .IN2(n533), .IN3(n527), .IN4(n517), .IN5(n800), 
        .Q(n799) );
  OA222X1 U751 ( .IN1(n528), .IN2(n542), .IN3(n523), .IN4(n516), .IN5(n530), 
        .IN6(n534), .Q(n800) );
  NAND3X0 U752 ( .IN1(N200), .IN2(n801), .IN3(n802), .QN(n530) );
  NAND3X0 U753 ( .IN1(n801), .IN2(n803), .IN3(n804), .QN(n516) );
  NAND3X0 U754 ( .IN1(n804), .IN2(n801), .IN3(n802), .QN(n528) );
  INVX0 U755 ( .INP(n574), .ZN(n527) );
  NOR3X0 U756 ( .IN1(n805), .IN2(n802), .IN3(n804), .QN(n574) );
  NAND2X0 U757 ( .IN1(N200), .IN2(N20), .QN(n804) );
  NAND3X0 U758 ( .IN1(n805), .IN2(n806), .IN3(n802), .QN(n533) );
  OA22X1 U759 ( .IN1(n525), .IN2(n537), .IN3(n521), .IN4(n536), .Q(n798) );
  NAND3X0 U760 ( .IN1(n803), .IN2(n806), .IN3(n805), .QN(n521) );
  NAND3X0 U761 ( .IN1(N200), .IN2(n803), .IN3(n805), .QN(n525) );
  INVX0 U762 ( .INP(n802), .ZN(n803) );
  NAND2X0 U763 ( .IN1(N68), .IN2(n712), .QN(n797) );
  INVX0 U764 ( .INP(n518), .ZN(n712) );
  NAND3X0 U765 ( .IN1(n805), .IN2(N200), .IN3(n802), .QN(n518) );
  NOR2X0 U766 ( .IN1(n779), .IN2(N190), .QN(n802) );
  INVX0 U767 ( .INP(n801), .ZN(n805) );
  NAND2X0 U768 ( .IN1(N179), .IN2(N20), .QN(n801) );
  NOR2X0 U769 ( .IN1(n558), .IN2(N33), .QN(n546) );
  AO21X1 U770 ( .IN1(N20), .IN2(n807), .IN3(n808), .Q(n558) );
  OR2X1 U771 ( .IN1(n780), .IN2(n715), .Q(n781) );
  INVX0 U772 ( .INP(n617), .ZN(n715) );
  NOR2X0 U773 ( .IN1(n548), .IN2(N20), .QN(n617) );
  INVX0 U774 ( .INP(n765), .ZN(n548) );
  NOR2X0 U775 ( .IN1(N33), .IN2(N13), .QN(n765) );
  AO21X1 U776 ( .IN1(n696), .IN2(n809), .IN3(n810), .Q(N4667) );
  MUX21X1 U777 ( .IN1(n811), .IN2(n812), .S(n623), .Q(n810) );
  NAND2X0 U778 ( .IN1(n796), .IN2(n563), .QN(n623) );
  NOR2X0 U779 ( .IN1(n809), .IN2(n674), .QN(n812) );
  NAND3X0 U780 ( .IN1(n519), .IN2(n517), .IN3(n813), .QN(n674) );
  INVX0 U781 ( .INP(n795), .ZN(n811) );
  INVX0 U782 ( .INP(n686), .ZN(n696) );
  NOR2X0 U783 ( .IN1(n649), .IN2(n738), .QN(n686) );
  INVX0 U784 ( .INP(n760), .ZN(n738) );
  NAND2X0 U785 ( .IN1(n814), .IN2(n742), .QN(n760) );
  NOR2X0 U786 ( .IN1(n815), .IN2(n816), .QN(n649) );
  INVX0 U787 ( .INP(N330), .ZN(n816) );
  MUX21X1 U788 ( .IN1(n817), .IN2(n818), .S(n742), .Q(n815) );
  MUX21X1 U789 ( .IN1(n819), .IN2(n820), .S(N179), .Q(n817) );
  OR4X1 U790 ( .IN1(n821), .IN2(n822), .IN3(n823), .IN4(n824), .Q(n820) );
  NAND4X0 U791 ( .IN1(n822), .IN2(n821), .IN3(n823), .IN4(n824), .QN(n819) );
  INVX0 U792 ( .INP(n695), .ZN(N4589) );
  OA22X1 U793 ( .IN1(n825), .IN2(n718), .IN3(n679), .IN4(n697), .Q(n695) );
  AOI22X1 U794 ( .IN1(n826), .IN2(n742), .IN3(N330), .IN4(n780), .QN(n697) );
  XNOR2X1 U795 ( .IN1(n827), .IN2(n828), .Q(n780) );
  NAND2X0 U796 ( .IN1(n718), .IN2(n829), .QN(n827) );
  XNOR2X1 U797 ( .IN1(n830), .IN2(n831), .Q(n679) );
  NOR2X0 U798 ( .IN1(n832), .IN2(n742), .QN(n831) );
  INVX0 U799 ( .INP(n718), .ZN(n742) );
  NOR2X0 U800 ( .IN1(n495), .IN2(n595), .QN(n718) );
  NAND4X0 U801 ( .IN1(N213), .IN2(N13), .IN3(n809), .IN4(n779), .QN(n595) );
  INVX0 U802 ( .INP(N343), .ZN(n495) );
  AO21X1 U803 ( .IN1(n650), .IN2(n814), .IN3(n739), .Q(N4145) );
  XOR2X1 U804 ( .IN1(keyinput22), .IN2(n833), .Q(n739) );
  OA21X1 U805 ( .IN1(n834), .IN2(n592), .IN3(n835), .Q(n833) );
  INVX0 U806 ( .INP(n836), .ZN(n592) );
  OA21X1 U807 ( .IN1(n837), .IN2(n838), .IN3(n839), .Q(n834) );
  INVX0 U808 ( .INP(n740), .ZN(n839) );
  AOI21X1 U809 ( .IN1(n746), .IN2(n743), .IN3(n741), .QN(n837) );
  INVX0 U810 ( .INP(n840), .ZN(n741) );
  NAND3X0 U811 ( .IN1(n841), .IN2(n842), .IN3(n843), .QN(n814) );
  NAND2X0 U812 ( .IN1(n723), .IN2(n844), .QN(n843) );
  AO21X1 U813 ( .IN1(n721), .IN2(n845), .IN3(n846), .Q(n844) );
  INVX0 U814 ( .INP(n719), .ZN(n846) );
  AO21X1 U815 ( .IN1(n830), .IN2(n826), .IN3(n847), .Q(n845) );
  INVX0 U816 ( .INP(n825), .ZN(n847) );
  INVX0 U817 ( .INP(n735), .ZN(n650) );
  NOR2X0 U818 ( .IN1(n735), .IN2(n818), .QN(N4028) );
  NAND4X0 U819 ( .IN1(n828), .IN2(n723), .IN3(n721), .IN4(n830), .QN(n818) );
  AND2X1 U820 ( .IN1(n848), .IN2(n825), .Q(n830) );
  NAND2X0 U821 ( .IN1(n849), .IN2(n850), .QN(n825) );
  MUX21X1 U822 ( .IN1(N179), .IN2(N169), .S(n822), .Q(n849) );
  NAND3X0 U823 ( .IN1(n851), .IN2(n852), .IN3(n832), .QN(n848) );
  INVX0 U824 ( .INP(n850), .ZN(n832) );
  AO221X1 U825 ( .IN1(n853), .IN2(N116), .IN3(n854), .IN4(N87), .IN5(n855), 
        .Q(n850) );
  MUX21X1 U826 ( .IN1(n856), .IN2(n857), .S(n534), .Q(n855) );
  NAND2X0 U827 ( .IN1(n858), .IN2(N190), .QN(n852) );
  XOR2X1 U828 ( .IN1(keyinput20), .IN2(n859), .Q(n851) );
  NOR2X0 U829 ( .IN1(n858), .IN2(n806), .QN(n859) );
  INVX0 U830 ( .INP(n822), .ZN(n858) );
  AO221X1 U831 ( .IN1(n860), .IN2(n861), .IN3(N264), .IN4(n862), .IN5(n863), 
        .Q(n822) );
  AO222X1 U832 ( .IN1(N250), .IN2(n864), .IN3(N257), .IN4(n865), .IN5(N294), 
        .IN6(N33), .Q(n861) );
  AND2X1 U833 ( .IN1(n866), .IN2(n719), .Q(n721) );
  NAND3X0 U834 ( .IN1(n867), .IN2(n722), .IN3(n868), .QN(n719) );
  MUX21X1 U835 ( .IN1(n869), .IN2(n823), .S(keyinput15), .Q(n868) );
  NAND2X0 U836 ( .IN1(n823), .IN2(n807), .QN(n869) );
  INVX0 U837 ( .INP(N169), .ZN(n807) );
  AO21X1 U838 ( .IN1(N169), .IN2(n823), .IN3(N179), .Q(n867) );
  AO221X1 U839 ( .IN1(N190), .IN2(n870), .IN3(N200), .IN4(n823), .IN5(n722), 
        .Q(n866) );
  AO221X1 U840 ( .IN1(n813), .IN2(n871), .IN3(n853), .IN4(N107), .IN5(n872), 
        .Q(n722) );
  OAI21X1 U841 ( .IN1(n531), .IN2(n873), .IN3(n874), .QN(n872) );
  MUX21X1 U842 ( .IN1(n875), .IN2(n876), .S(n523), .Q(n874) );
  OA21X1 U843 ( .IN1(n534), .IN2(n877), .IN3(n878), .Q(n875) );
  INVX0 U844 ( .INP(N107), .ZN(n534) );
  XNOR2X1 U845 ( .IN1(keyinput15), .IN2(n823), .Q(n870) );
  AO221X1 U846 ( .IN1(n860), .IN2(n879), .IN3(N257), .IN4(n862), .IN5(n863), 
        .Q(n823) );
  AO222X1 U847 ( .IN1(N244), .IN2(n864), .IN3(N250), .IN4(n865), .IN5(N283), 
        .IN6(N33), .Q(n879) );
  AND3X1 U848 ( .IN1(n841), .IN2(n842), .IN3(n880), .Q(n723) );
  NAND2X0 U849 ( .IN1(n881), .IN2(n882), .QN(n880) );
  XOR2X1 U850 ( .IN1(n725), .IN2(keyinput10), .Q(n882) );
  MUX21X1 U851 ( .IN1(n883), .IN2(n806), .S(n824), .Q(n881) );
  NAND3X0 U852 ( .IN1(N179), .IN2(n725), .IN3(n884), .QN(n842) );
  INVX0 U853 ( .INP(n824), .ZN(n884) );
  NAND3X0 U854 ( .IN1(n725), .IN2(n824), .IN3(N169), .QN(n841) );
  AO21X1 U855 ( .IN1(n885), .IN2(N274), .IN3(n886), .Q(n824) );
  MUX21X1 U856 ( .IN1(n887), .IN2(n888), .S(n860), .Q(n886) );
  AO222X1 U857 ( .IN1(N238), .IN2(n864), .IN3(N244), .IN4(n865), .IN5(N116), 
        .IN6(N33), .Q(n888) );
  NOR2X0 U858 ( .IN1(n885), .IN2(n889), .QN(n887) );
  NAND4X0 U859 ( .IN1(n890), .IN2(n891), .IN3(n892), .IN4(n893), .QN(n725) );
  NAND3X0 U860 ( .IN1(n894), .IN2(n895), .IN3(N97), .QN(n893) );
  NAND2X0 U861 ( .IN1(N68), .IN2(n854), .QN(n892) );
  NAND2X0 U862 ( .IN1(n871), .IN2(N107), .QN(n891) );
  MUX21X1 U863 ( .IN1(n896), .IN2(n876), .S(n517), .Q(n890) );
  NOR2X0 U864 ( .IN1(n871), .IN2(n856), .QN(n896) );
  INVX0 U865 ( .INP(n878), .ZN(n856) );
  AOI21X1 U866 ( .IN1(n897), .IN2(n898), .IN3(n826), .QN(n828) );
  AND2X1 U867 ( .IN1(n899), .IN2(n829), .Q(n826) );
  MUX21X1 U868 ( .IN1(N179), .IN2(N169), .S(n821), .Q(n899) );
  INVX0 U869 ( .INP(n829), .ZN(n898) );
  NAND3X0 U870 ( .IN1(n900), .IN2(n901), .IN3(n902), .QN(n829) );
  OA22X1 U871 ( .IN1(n522), .IN2(n903), .IN3(n523), .IN4(n873), .Q(n902) );
  INVX0 U872 ( .INP(N97), .ZN(n523) );
  INVX0 U873 ( .INP(N283), .ZN(n522) );
  XOR2X1 U874 ( .IN1(keyinput4), .IN2(n904), .Q(n901) );
  NOR2X0 U875 ( .IN1(n519), .IN2(n878), .QN(n904) );
  NAND3X0 U876 ( .IN1(n905), .IN2(n876), .IN3(n906), .QN(n878) );
  NAND2X0 U877 ( .IN1(n907), .IN2(n809), .QN(n905) );
  XNOR2X1 U878 ( .IN1(keyinput0), .IN2(n566), .Q(n907) );
  MUX21X1 U879 ( .IN1(n877), .IN2(n876), .S(n519), .Q(n900) );
  INVX0 U880 ( .INP(N116), .ZN(n519) );
  MUX21X1 U881 ( .IN1(n883), .IN2(n806), .S(n821), .Q(n897) );
  AO221X1 U882 ( .IN1(n860), .IN2(n908), .IN3(N270), .IN4(n862), .IN5(n863), 
        .Q(n821) );
  AND3X1 U883 ( .IN1(N274), .IN2(n563), .IN3(n885), .Q(n863) );
  AOI21X1 U884 ( .IN1(n885), .IN2(n563), .IN3(n860), .QN(n862) );
  NOR2X0 U885 ( .IN1(n672), .IN2(N1), .QN(n885) );
  AO222X1 U886 ( .IN1(N257), .IN2(n864), .IN3(N264), .IN4(n865), .IN5(N303), 
        .IN6(N33), .Q(n908) );
  NAND4X0 U887 ( .IN1(n748), .IN2(n772), .IN3(n836), .IN4(n746), .QN(n735) );
  OA21X1 U888 ( .IN1(n909), .IN2(n747), .IN3(n840), .Q(n746) );
  NAND2X0 U889 ( .IN1(n910), .IN2(n747), .QN(n840) );
  MUX21X1 U890 ( .IN1(N169), .IN2(N179), .S(n911), .Q(n910) );
  AO221X1 U891 ( .IN1(n853), .IN2(N77), .IN3(n854), .IN4(N50), .IN5(n912), .Q(
        n747) );
  MUX21X1 U892 ( .IN1(n913), .IN2(n857), .S(n513), .Q(n912) );
  NAND2X0 U893 ( .IN1(n876), .IN2(n877), .QN(n857) );
  MUX21X1 U894 ( .IN1(N200), .IN2(N190), .S(n911), .Q(n909) );
  AOI221X1 U895 ( .IN1(n860), .IN2(n914), .IN3(N238), .IN4(n915), .IN5(n916), 
        .QN(n911) );
  AO222X1 U896 ( .IN1(N226), .IN2(n864), .IN3(N232), .IN4(n865), .IN5(N97), 
        .IN6(N33), .Q(n914) );
  OA21X1 U897 ( .IN1(n917), .IN2(n594), .IN3(n835), .Q(n836) );
  NAND2X0 U898 ( .IN1(n918), .IN2(n594), .QN(n835) );
  MUX21X1 U899 ( .IN1(N169), .IN2(N179), .S(n919), .Q(n918) );
  NAND4X0 U900 ( .IN1(n920), .IN2(n921), .IN3(n922), .IN4(n923), .QN(n594) );
  NAND3X0 U901 ( .IN1(n894), .IN2(n895), .IN3(N58), .QN(n923) );
  NAND2X0 U902 ( .IN1(n854), .IN2(N150), .QN(n922) );
  NAND2X0 U903 ( .IN1(n871), .IN2(N68), .QN(n921) );
  MUX21X1 U904 ( .IN1(n924), .IN2(n876), .S(n537), .Q(n920) );
  MUX21X1 U905 ( .IN1(N200), .IN2(N190), .S(n919), .Q(n917) );
  AOI221X1 U906 ( .IN1(n860), .IN2(n925), .IN3(n915), .IN4(N226), .IN5(n916), 
        .QN(n919) );
  AO222X1 U907 ( .IN1(N222), .IN2(n864), .IN3(N223), .IN4(n865), .IN5(N77), 
        .IN6(N33), .Q(n925) );
  AOI21X1 U908 ( .IN1(n926), .IN2(n927), .IN3(n743), .QN(n772) );
  AND2X1 U909 ( .IN1(n928), .IN2(n773), .Q(n743) );
  INVX0 U910 ( .INP(n927), .ZN(n773) );
  MUX21X1 U911 ( .IN1(N169), .IN2(N179), .S(n929), .Q(n928) );
  OA221X1 U912 ( .IN1(n903), .IN2(n517), .IN3(n873), .IN4(n536), .IN5(n930), 
        .Q(n927) );
  MUX21X1 U913 ( .IN1(n924), .IN2(n876), .S(n531), .Q(n930) );
  INVX0 U914 ( .INP(N77), .ZN(n531) );
  NOR2X0 U915 ( .IN1(n913), .IN2(n871), .QN(n924) );
  MUX21X1 U916 ( .IN1(n806), .IN2(n883), .S(n929), .Q(n926) );
  AOI221X1 U917 ( .IN1(n860), .IN2(n931), .IN3(N244), .IN4(n915), .IN5(n916), 
        .QN(n929) );
  AO222X1 U918 ( .IN1(n864), .IN2(N232), .IN3(N238), .IN4(n865), .IN5(N107), 
        .IN6(N33), .Q(n931) );
  INVX0 U919 ( .INP(n838), .ZN(n748) );
  AO21X1 U920 ( .IN1(n932), .IN2(n750), .IN3(n740), .Q(n838) );
  NOR2X0 U921 ( .IN1(n933), .IN2(n750), .QN(n740) );
  INVX0 U922 ( .INP(n934), .ZN(n933) );
  MUX21X1 U923 ( .IN1(N169), .IN2(N179), .S(n935), .Q(n934) );
  OA221X1 U924 ( .IN1(n936), .IN2(n513), .IN3(n542), .IN4(n873), .IN5(n937), 
        .Q(n750) );
  MUX21X1 U925 ( .IN1(n938), .IN2(n939), .S(n536), .Q(n937) );
  OA21X1 U926 ( .IN1(N68), .IN2(n877), .IN3(n876), .Q(n939) );
  NAND2X0 U927 ( .IN1(n940), .IN2(N13), .QN(n876) );
  INVX0 U928 ( .INP(n913), .ZN(n938) );
  NOR2X0 U929 ( .IN1(n894), .IN2(n940), .QN(n913) );
  NOR2X0 U930 ( .IN1(n779), .IN2(N1), .QN(n940) );
  INVX0 U931 ( .INP(n854), .ZN(n873) );
  NOR2X0 U932 ( .IN1(n895), .IN2(n906), .QN(n854) );
  NAND2X0 U933 ( .IN1(n941), .IN2(n779), .QN(n895) );
  INVX0 U934 ( .INP(N159), .ZN(n542) );
  OA21X1 U935 ( .IN1(n536), .IN2(n877), .IN3(n903), .Q(n936) );
  INVX0 U936 ( .INP(n853), .ZN(n903) );
  NOR2X0 U937 ( .IN1(n941), .IN2(n906), .QN(n853) );
  NAND2X0 U938 ( .IN1(N33), .IN2(n779), .QN(n941) );
  INVX0 U939 ( .INP(n871), .ZN(n877) );
  NOR2X0 U940 ( .IN1(n779), .IN2(n906), .QN(n871) );
  INVX0 U941 ( .INP(n894), .ZN(n906) );
  NAND2X0 U942 ( .IN1(n808), .IN2(n942), .QN(n894) );
  NAND3X0 U943 ( .IN1(N20), .IN2(N1), .IN3(N33), .QN(n942) );
  INVX0 U944 ( .INP(N20), .ZN(n779) );
  MUX21X1 U945 ( .IN1(n806), .IN2(n883), .S(n935), .Q(n932) );
  AOI221X1 U946 ( .IN1(n943), .IN2(n860), .IN3(n915), .IN4(N232), .IN5(n916), 
        .QN(n935) );
  AND3X1 U947 ( .IN1(n944), .IN2(n809), .IN3(N274), .Q(n916) );
  AOI21X1 U948 ( .IN1(n809), .IN2(n944), .IN3(n860), .QN(n915) );
  NAND2X0 U949 ( .IN1(n672), .IN2(n563), .QN(n944) );
  INVX0 U950 ( .INP(N45), .ZN(n672) );
  OA21X1 U951 ( .IN1(n563), .IN2(n566), .IN3(n945), .Q(n860) );
  INVX0 U952 ( .INP(N33), .ZN(n566) );
  INVX0 U953 ( .INP(N41), .ZN(n563) );
  XOR2X1 U954 ( .IN1(n946), .IN2(keyinput7), .Q(n943) );
  AO221X1 U955 ( .IN1(N226), .IN2(n865), .IN3(N87), .IN4(N33), .IN5(n947), .Q(
        n946) );
  XOR2X1 U956 ( .IN1(keyinput2), .IN2(n948), .Q(n947) );
  AND2X1 U957 ( .IN1(n864), .IN2(N223), .Q(n948) );
  NOR2X0 U958 ( .IN1(n864), .IN2(N33), .QN(n865) );
  NOR2X0 U959 ( .IN1(N349), .IN2(N33), .QN(n864) );
  INVX0 U960 ( .INP(N190), .ZN(n883) );
  INVX0 U961 ( .INP(N200), .ZN(n806) );
  MUX21X1 U962 ( .IN1(n949), .IN2(n950), .S(n613), .Q(N3987) );
  XNOR3X1 U963 ( .IN1(N97), .IN2(n951), .IN3(n517), .Q(n613) );
  NOR2X0 U964 ( .IN1(keyinput8), .IN2(n952), .QN(n951) );
  XNOR2X1 U965 ( .IN1(N116), .IN2(N107), .Q(n952) );
  OR2X1 U966 ( .IN1(n794), .IN2(keyinput21), .Q(n950) );
  INVX0 U967 ( .INP(n949), .ZN(n794) );
  AO21X1 U968 ( .IN1(n953), .IN2(n954), .IN3(n955), .Q(n949) );
  MUX21X1 U969 ( .IN1(n956), .IN2(n957), .S(n536), .Q(n955) );
  XNOR2X1 U970 ( .IN1(n537), .IN2(n954), .Q(n957) );
  NOR2X0 U971 ( .IN1(N50), .IN2(n954), .QN(n956) );
  AOI21X1 U972 ( .IN1(N77), .IN2(n513), .IN3(n958), .QN(n954) );
  XOR2X1 U973 ( .IN1(keyinput5), .IN2(n959), .Q(n958) );
  NOR2X0 U974 ( .IN1(N77), .IN2(n513), .QN(n959) );
  XOR2X1 U975 ( .IN1(n713), .IN2(n673), .Q(N3833) );
  XNOR3X1 U976 ( .IN1(N232), .IN2(N226), .IN3(n960), .Q(n673) );
  XNOR2X1 U977 ( .IN1(N238), .IN2(N244), .Q(n960) );
  XNOR3X1 U978 ( .IN1(N257), .IN2(n889), .IN3(n961), .Q(n713) );
  XNOR2X1 U979 ( .IN1(N270), .IN2(N264), .Q(n961) );
  INVX0 U980 ( .INP(N250), .ZN(n889) );
  OA21X1 U981 ( .IN1(n795), .IN2(n731), .IN3(n962), .Q(N3195) );
  MUX21X1 U982 ( .IN1(n963), .IN2(n964), .S(n796), .Q(n962) );
  AND2X1 U983 ( .IN1(N20), .IN2(n726), .Q(n796) );
  NOR2X0 U984 ( .IN1(n809), .IN2(N13), .QN(n726) );
  INVX0 U985 ( .INP(N1), .ZN(n809) );
  OAI21X1 U986 ( .IN1(N257), .IN2(N264), .IN3(N250), .QN(n964) );
  NAND2X0 U987 ( .IN1(n965), .IN2(n731), .QN(n963) );
  NAND4X0 U988 ( .IN1(n966), .IN2(n967), .IN3(n968), .IN4(n969), .QN(n965) );
  AOI221X1 U989 ( .IN1(N68), .IN2(N238), .IN3(N50), .IN4(N226), .IN5(n970), 
        .QN(n969) );
  AO22X1 U990 ( .IN1(N107), .IN2(N264), .IN3(N116), .IN4(N270), .Q(n970) );
  AOI22X1 U991 ( .IN1(N77), .IN2(N244), .IN3(N87), .IN4(N250), .QN(n968) );
  NAND2X0 U992 ( .IN1(N257), .IN2(N97), .QN(n967) );
  XOR2X1 U993 ( .IN1(n971), .IN2(keyinput1), .Q(n966) );
  NAND2X0 U994 ( .IN1(N232), .IN2(N58), .QN(n971) );
  NAND2X0 U995 ( .IN1(n945), .IN2(N20), .QN(n731) );
  INVX0 U996 ( .INP(n808), .ZN(n945) );
  NAND2X0 U997 ( .IN1(N13), .IN2(N1), .QN(n808) );
  OA21X1 U998 ( .IN1(n513), .IN2(n537), .IN3(n756), .Q(n795) );
  INVX0 U999 ( .INP(n953), .ZN(n756) );
  NOR2X0 U1000 ( .IN1(n536), .IN2(n537), .QN(n953) );
  INVX0 U1001 ( .INP(N58), .ZN(n536) );
  INVX0 U1002 ( .INP(N50), .ZN(n537) );
  INVX0 U1003 ( .INP(N68), .ZN(n513) );
  NOR4X0 U1004 ( .IN1(N77), .IN2(N68), .IN3(N58), .IN4(N50), .QN(N1713) );
  OR2X1 U1005 ( .IN1(n517), .IN2(n813), .Q(N1947) );
  NOR2X0 U1006 ( .IN1(N107), .IN2(N97), .QN(n813) );
  INVX0 U1007 ( .INP(N87), .ZN(n517) );
endmodule

