
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563;

  XNOR2X1 U331 ( .IN1(keyinput62), .IN2(n303), .Q(G1348) );
  OA22X1 U332 ( .IN1(n304), .IN2(n305), .IN3(G25), .IN4(n306), .Q(n303) );
  AND2X1 U333 ( .IN1(n307), .IN2(n304), .Q(n306) );
  OA21X1 U334 ( .IN1(n308), .IN2(n309), .IN3(n310), .Q(n304) );
  XNOR3X1 U335 ( .IN1(keyinput40), .IN2(G31), .IN3(n311), .Q(G1354) );
  NAND2X0 U336 ( .IN1(n312), .IN2(n313), .QN(n311) );
  XNOR2X1 U337 ( .IN1(n314), .IN2(n315), .Q(G1352) );
  NAND2X0 U338 ( .IN1(n312), .IN2(n310), .QN(n314) );
  OA21X1 U339 ( .IN1(G28), .IN2(n316), .IN3(n317), .Q(G1351) );
  XOR2X1 U340 ( .IN1(keyinput55), .IN2(n318), .Q(n317) );
  AND2X1 U341 ( .IN1(G28), .IN2(n316), .Q(n318) );
  XOR2X1 U342 ( .IN1(n319), .IN2(keyinput39), .Q(n316) );
  NAND2X0 U343 ( .IN1(n307), .IN2(n320), .QN(n319) );
  OA21X1 U344 ( .IN1(G26), .IN2(n321), .IN3(n322), .Q(G1349) );
  XOR2X1 U345 ( .IN1(keyinput53), .IN2(n323), .Q(n322) );
  AND2X1 U346 ( .IN1(n321), .IN2(G26), .Q(n323) );
  NAND2X0 U347 ( .IN1(n307), .IN2(n324), .QN(n321) );
  INVX0 U348 ( .INP(n308), .ZN(n307) );
  AOI21X1 U349 ( .IN1(n325), .IN2(G24), .IN3(n326), .QN(G1347) );
  AND3X1 U350 ( .IN1(n325), .IN2(n320), .IN3(n327), .Q(n326) );
  XNOR2X1 U351 ( .IN1(n328), .IN2(keyinput42), .Q(n325) );
  NAND3X0 U352 ( .IN1(G24), .IN2(n320), .IN3(n327), .QN(n328) );
  XOR3X1 U353 ( .IN1(keyinput38), .IN2(G23), .IN3(n329), .Q(G1346) );
  NAND2X0 U354 ( .IN1(n327), .IN2(n313), .QN(n329) );
  XNOR2X1 U355 ( .IN1(G22), .IN2(n330), .Q(G1345) );
  NOR2X0 U356 ( .IN1(n331), .IN2(n332), .QN(n330) );
  OA21X1 U357 ( .IN1(n333), .IN2(n334), .IN3(n335), .Q(G1344) );
  XOR2X1 U358 ( .IN1(n336), .IN2(keyinput52), .Q(n335) );
  NAND3X0 U359 ( .IN1(n310), .IN2(n334), .IN3(n327), .QN(n336) );
  INVX0 U360 ( .INP(n332), .ZN(n327) );
  NOR2X0 U361 ( .IN1(n305), .IN2(n332), .QN(n333) );
  NAND4X0 U362 ( .IN1(n337), .IN2(n338), .IN3(n339), .IN4(n340), .QN(n332) );
  NOR2X0 U363 ( .IN1(n341), .IN2(n342), .QN(n340) );
  OA21X1 U364 ( .IN1(n343), .IN2(n344), .IN3(n345), .Q(G1342) );
  XOR2X1 U365 ( .IN1(n346), .IN2(keyinput50), .Q(n345) );
  NAND2X0 U366 ( .IN1(n343), .IN2(n344), .QN(n346) );
  INVX0 U367 ( .INP(G19), .ZN(n344) );
  XOR2X1 U368 ( .IN1(n347), .IN2(keyinput37), .Q(n343) );
  NAND2X0 U369 ( .IN1(n348), .IN2(n313), .QN(n347) );
  XNOR2X1 U370 ( .IN1(G18), .IN2(n349), .Q(G1341) );
  NOR2X0 U371 ( .IN1(n331), .IN2(n350), .QN(n349) );
  MUX21X1 U372 ( .IN1(n351), .IN2(n352), .S(G17), .Q(G1340) );
  NOR2X0 U373 ( .IN1(n305), .IN2(n350), .QN(n352) );
  NAND2X0 U374 ( .IN1(n348), .IN2(n310), .QN(n351) );
  INVX0 U375 ( .INP(n350), .ZN(n348) );
  NOR2X0 U376 ( .IN1(n353), .IN2(n354), .QN(G1338) );
  XOR2X1 U377 ( .IN1(keyinput49), .IN2(n355), .Q(n354) );
  NOR2X0 U378 ( .IN1(G15), .IN2(n356), .QN(n355) );
  XOR2X1 U379 ( .IN1(n357), .IN2(keyinput48), .Q(n353) );
  NAND2X0 U380 ( .IN1(G15), .IN2(n356), .QN(n357) );
  NAND2X0 U381 ( .IN1(n358), .IN2(n342), .QN(n356) );
  XNOR2X1 U382 ( .IN1(n359), .IN2(n360), .Q(G1337) );
  NAND2X0 U383 ( .IN1(n358), .IN2(n341), .QN(n359) );
  OA21X1 U384 ( .IN1(G13), .IN2(n361), .IN3(n362), .Q(G1336) );
  XOR2X1 U385 ( .IN1(keyinput47), .IN2(n363), .Q(n362) );
  AND2X1 U386 ( .IN1(n361), .IN2(G13), .Q(n363) );
  NAND2X0 U387 ( .IN1(n358), .IN2(n338), .QN(n361) );
  XNOR2X1 U388 ( .IN1(G12), .IN2(n364), .Q(G1335) );
  NOR2X0 U389 ( .IN1(n365), .IN2(n366), .QN(n364) );
  NOR2X0 U390 ( .IN1(n367), .IN2(n368), .QN(G1334) );
  XOR2X1 U391 ( .IN1(keyinput46), .IN2(n369), .Q(n368) );
  NOR2X0 U392 ( .IN1(n370), .IN2(n371), .QN(n369) );
  NOR3X0 U393 ( .IN1(n366), .IN2(n370), .IN3(n372), .QN(n367) );
  NOR3X0 U394 ( .IN1(n371), .IN2(n372), .IN3(n366), .QN(n370) );
  NOR2X0 U395 ( .IN1(n373), .IN2(n374), .QN(G1333) );
  XOR2X1 U396 ( .IN1(keyinput45), .IN2(n375), .Q(n374) );
  NOR2X0 U397 ( .IN1(n376), .IN2(n377), .QN(n375) );
  NOR3X0 U398 ( .IN1(n366), .IN2(n376), .IN3(n378), .QN(n373) );
  NOR3X0 U399 ( .IN1(n377), .IN2(n378), .IN3(n366), .QN(n376) );
  OA21X1 U400 ( .IN1(n379), .IN2(n380), .IN3(n381), .Q(G1332) );
  XOR2X1 U401 ( .IN1(n382), .IN2(keyinput44), .Q(n381) );
  OR3X1 U402 ( .IN1(n383), .IN2(G9), .IN3(n366), .Q(n382) );
  INVX0 U403 ( .INP(G9), .ZN(n380) );
  NOR2X0 U404 ( .IN1(n383), .IN2(n366), .QN(n379) );
  NAND4X0 U405 ( .IN1(n384), .IN2(n313), .IN3(n305), .IN4(n385), .QN(n366) );
  NOR2X0 U406 ( .IN1(n320), .IN2(n331), .QN(n385) );
  XNOR2X1 U407 ( .IN1(G8), .IN2(n386), .Q(G1331) );
  NOR2X0 U408 ( .IN1(n365), .IN2(n387), .QN(n386) );
  XNOR2X1 U409 ( .IN1(G7), .IN2(n388), .Q(G1330) );
  NOR2X0 U410 ( .IN1(n372), .IN2(n387), .QN(n388) );
  XNOR2X1 U411 ( .IN1(G6), .IN2(n389), .Q(G1329) );
  NOR2X0 U412 ( .IN1(n378), .IN2(n387), .QN(n389) );
  XNOR2X1 U413 ( .IN1(G5), .IN2(n390), .Q(G1328) );
  NOR2X0 U414 ( .IN1(n383), .IN2(n387), .QN(n390) );
  NAND4X0 U415 ( .IN1(n320), .IN2(n384), .IN3(n331), .IN4(n391), .QN(n387) );
  NOR2X0 U416 ( .IN1(n313), .IN2(n305), .QN(n391) );
  XOR2X1 U417 ( .IN1(n392), .IN2(G4), .Q(G1327) );
  NAND2X0 U418 ( .IN1(n393), .IN2(n339), .QN(n392) );
  OA21X1 U419 ( .IN1(n394), .IN2(n395), .IN3(n396), .Q(G1325) );
  XOR2X1 U420 ( .IN1(n397), .IN2(keyinput43), .Q(n396) );
  NAND2X0 U421 ( .IN1(n398), .IN2(n399), .QN(n397) );
  INVX0 U422 ( .INP(n395), .ZN(n398) );
  XNOR2X1 U423 ( .IN1(n400), .IN2(keyinput41), .Q(n395) );
  NAND2X0 U424 ( .IN1(n399), .IN2(G2), .QN(n400) );
  NOR2X0 U425 ( .IN1(n401), .IN2(n378), .QN(n399) );
  XNOR2X1 U426 ( .IN1(n402), .IN2(n403), .Q(G1324) );
  NAND2X0 U427 ( .IN1(n393), .IN2(n338), .QN(n402) );
  XNOR2X1 U428 ( .IN1(keyinput59), .IN2(n404), .Q(G1350) );
  NOR2X0 U429 ( .IN1(n405), .IN2(n406), .QN(n404) );
  XOR2X1 U430 ( .IN1(n407), .IN2(keyinput54), .Q(n406) );
  OR3X1 U431 ( .IN1(n408), .IN2(G27), .IN3(n308), .Q(n407) );
  OA21X1 U432 ( .IN1(n408), .IN2(n308), .IN3(G27), .Q(n405) );
  NAND3X0 U433 ( .IN1(n409), .IN2(n341), .IN3(n383), .QN(n308) );
  XOR3X1 U434 ( .IN1(keyinput60), .IN2(G32), .IN3(n410), .Q(G1355) );
  NAND2X0 U435 ( .IN1(n312), .IN2(n320), .QN(n410) );
  XOR2X1 U436 ( .IN1(keyinput63), .IN2(n411), .Q(G1353) );
  OA21X1 U437 ( .IN1(G30), .IN2(n412), .IN3(n413), .Q(n411) );
  XOR2X1 U438 ( .IN1(n414), .IN2(n415), .Q(n413) );
  NOR2X0 U439 ( .IN1(keyinput56), .IN2(n416), .QN(n415) );
  NAND2X0 U440 ( .IN1(n312), .IN2(n324), .QN(n414) );
  AND4X1 U441 ( .IN1(n372), .IN2(n417), .IN3(n383), .IN4(n337), .Q(n312) );
  INVX0 U442 ( .INP(keyinput56), .ZN(n412) );
  XOR2X1 U443 ( .IN1(keyinput58), .IN2(n418), .Q(G1343) );
  OA21X1 U444 ( .IN1(G20), .IN2(n419), .IN3(n420), .Q(n418) );
  XOR2X1 U445 ( .IN1(n421), .IN2(n422), .Q(n420) );
  NOR2X0 U446 ( .IN1(n423), .IN2(n350), .QN(n422) );
  NAND3X0 U447 ( .IN1(n409), .IN2(n338), .IN3(n378), .QN(n350) );
  AND3X1 U448 ( .IN1(n342), .IN2(n337), .IN3(n365), .Q(n409) );
  NAND2X0 U449 ( .IN1(n424), .IN2(n425), .QN(n337) );
  OR3X1 U450 ( .IN1(n310), .IN2(n426), .IN3(n313), .Q(n425) );
  INVX0 U451 ( .INP(n305), .ZN(n310) );
  OR3X1 U452 ( .IN1(n324), .IN2(n427), .IN3(n320), .Q(n424) );
  NAND2X0 U453 ( .IN1(G20), .IN2(n419), .QN(n421) );
  INVX0 U454 ( .INP(keyinput51), .ZN(n419) );
  XNOR2X1 U455 ( .IN1(keyinput57), .IN2(n428), .Q(G1339) );
  OA22X1 U456 ( .IN1(n429), .IN2(n365), .IN3(G16), .IN4(n430), .Q(n428) );
  NOR2X0 U457 ( .IN1(n431), .IN2(n432), .QN(n430) );
  INVX0 U458 ( .INP(n432), .ZN(n429) );
  AO21X1 U459 ( .IN1(n358), .IN2(G16), .IN3(n365), .Q(n432) );
  INVX0 U460 ( .INP(n431), .ZN(n358) );
  NAND4X0 U461 ( .IN1(n433), .IN2(n426), .IN3(n305), .IN4(n384), .QN(n431) );
  NOR2X0 U462 ( .IN1(n331), .IN2(n423), .QN(n426) );
  XNOR2X1 U463 ( .IN1(n408), .IN2(keyinput35), .Q(n433) );
  XOR2X1 U464 ( .IN1(keyinput61), .IN2(n434), .Q(G1326) );
  OA22X1 U465 ( .IN1(n435), .IN2(n372), .IN3(G3), .IN4(n436), .Q(n434) );
  NOR2X0 U466 ( .IN1(n401), .IN2(n437), .QN(n436) );
  INVX0 U467 ( .INP(n437), .ZN(n435) );
  AO21X1 U468 ( .IN1(n393), .IN2(G3), .IN3(n372), .Q(n437) );
  INVX0 U469 ( .INP(n401), .ZN(n393) );
  NAND4X0 U470 ( .IN1(n438), .IN2(n427), .IN3(n423), .IN4(n384), .QN(n401) );
  AO222X1 U471 ( .IN1(n439), .IN2(n372), .IN3(n440), .IN4(n378), .IN5(
        keyinput36), .IN6(n441), .Q(n384) );
  NAND3X0 U472 ( .IN1(n365), .IN2(n383), .IN3(n378), .QN(n441) );
  INVX0 U473 ( .INP(n338), .ZN(n383) );
  NOR2X0 U474 ( .IN1(n442), .IN2(n339), .QN(n440) );
  OA21X1 U475 ( .IN1(keyinput36), .IN2(n338), .IN3(n342), .Q(n442) );
  INVX0 U476 ( .INP(n342), .ZN(n372) );
  XNOR3X1 U477 ( .IN1(n443), .IN2(n444), .IN3(n445), .Q(n342) );
  XNOR2X1 U478 ( .IN1(n446), .IN2(n447), .Q(n445) );
  OA21X1 U479 ( .IN1(G15), .IN2(n371), .IN3(n448), .Q(n447) );
  XOR2X1 U480 ( .IN1(keyinput9), .IN2(n449), .Q(n448) );
  AND2X1 U481 ( .IN1(n371), .IN2(G15), .Q(n449) );
  INVX0 U482 ( .INP(G11), .ZN(n371) );
  XNOR3X1 U483 ( .IN1(G7), .IN2(G3), .IN3(n450), .Q(n444) );
  NAND2X0 U484 ( .IN1(G35), .IN2(G41), .QN(n450) );
  NOR2X0 U485 ( .IN1(n417), .IN2(n338), .QN(n439) );
  AO21X1 U486 ( .IN1(n451), .IN2(n452), .IN3(n453), .Q(n338) );
  XOR2X1 U487 ( .IN1(keyinput31), .IN2(n454), .Q(n453) );
  NOR2X0 U488 ( .IN1(n451), .IN2(n452), .QN(n454) );
  XNOR3X1 U489 ( .IN1(G9), .IN2(n455), .IN3(G13), .Q(n452) );
  OA21X1 U490 ( .IN1(G5), .IN2(n403), .IN3(n456), .Q(n455) );
  XOR2X1 U491 ( .IN1(n457), .IN2(keyinput7), .Q(n456) );
  NAND2X0 U492 ( .IN1(G5), .IN2(n403), .QN(n457) );
  INVX0 U493 ( .INP(G1), .ZN(n403) );
  XOR3X1 U494 ( .IN1(keyinput25), .IN2(keyinput0), .IN3(n458), .Q(n451) );
  XOR2X1 U495 ( .IN1(n459), .IN2(n460), .Q(n458) );
  OA21X1 U496 ( .IN1(n461), .IN2(n443), .IN3(n462), .Q(n460) );
  XOR2X1 U497 ( .IN1(n463), .IN2(keyinput22), .Q(n462) );
  NAND2X0 U498 ( .IN1(n461), .IN2(n443), .QN(n463) );
  XNOR3X1 U499 ( .IN1(G18), .IN2(G17), .IN3(n464), .Q(n443) );
  XNOR3X1 U500 ( .IN1(keyinput18), .IN2(G20), .IN3(G19), .Q(n464) );
  NAND2X0 U501 ( .IN1(G41), .IN2(G33), .QN(n459) );
  NOR2X0 U502 ( .IN1(n378), .IN2(n365), .QN(n417) );
  INVX0 U503 ( .INP(n339), .ZN(n365) );
  XNOR3X1 U504 ( .IN1(n465), .IN2(n466), .IN3(n467), .Q(n339) );
  XNOR2X1 U505 ( .IN1(G4), .IN2(G8), .Q(n467) );
  OA21X1 U506 ( .IN1(G16), .IN2(n468), .IN3(n469), .Q(n466) );
  XOR2X1 U507 ( .IN1(n470), .IN2(keyinput10), .Q(n469) );
  NAND2X0 U508 ( .IN1(G16), .IN2(n468), .QN(n470) );
  INVX0 U509 ( .INP(G12), .ZN(n468) );
  OA21X1 U510 ( .IN1(n471), .IN2(n472), .IN3(n473), .Q(n465) );
  XOR2X1 U511 ( .IN1(keyinput29), .IN2(n474), .Q(n473) );
  NOR2X0 U512 ( .IN1(n471), .IN2(n475), .QN(n474) );
  NOR2X0 U513 ( .IN1(n475), .IN2(n472), .QN(n471) );
  XOR2X1 U514 ( .IN1(n476), .IN2(n461), .Q(n472) );
  XNOR3X1 U515 ( .IN1(G22), .IN2(n334), .IN3(n477), .Q(n461) );
  XNOR2X1 U516 ( .IN1(G23), .IN2(G24), .Q(n477) );
  NAND2X0 U517 ( .IN1(G36), .IN2(G41), .QN(n475) );
  INVX0 U518 ( .INP(n341), .ZN(n378) );
  XNOR2X1 U519 ( .IN1(n478), .IN2(keyinput33), .Q(n341) );
  NAND2X0 U520 ( .IN1(n479), .IN2(n480), .QN(n478) );
  NAND3X0 U521 ( .IN1(n481), .IN2(n482), .IN3(n483), .QN(n480) );
  XNOR2X1 U522 ( .IN1(keyinput30), .IN2(n484), .Q(n479) );
  AOI21X1 U523 ( .IN1(n481), .IN2(n482), .IN3(n483), .QN(n484) );
  XNOR3X1 U524 ( .IN1(n446), .IN2(n485), .IN3(n476), .Q(n483) );
  AO21X1 U525 ( .IN1(n486), .IN2(n487), .IN3(n488), .Q(n476) );
  XOR2X1 U526 ( .IN1(n489), .IN2(keyinput16), .Q(n488) );
  OR2X1 U527 ( .IN1(n487), .IN2(n486), .Q(n489) );
  AO21X1 U528 ( .IN1(n315), .IN2(n416), .IN3(n490), .Q(n487) );
  XOR2X1 U529 ( .IN1(keyinput3), .IN2(n491), .Q(n490) );
  NOR2X0 U530 ( .IN1(n416), .IN2(n315), .QN(n491) );
  XOR2X1 U531 ( .IN1(G31), .IN2(G32), .Q(n486) );
  XNOR2X1 U532 ( .IN1(n492), .IN2(keyinput26), .Q(n485) );
  NAND2X0 U533 ( .IN1(G34), .IN2(G41), .QN(n492) );
  XNOR3X1 U534 ( .IN1(G26), .IN2(G25), .IN3(n493), .Q(n446) );
  XNOR3X1 U535 ( .IN1(keyinput13), .IN2(G28), .IN3(G27), .Q(n493) );
  NAND2X0 U536 ( .IN1(n494), .IN2(n495), .QN(n482) );
  NAND2X0 U537 ( .IN1(n496), .IN2(n495), .QN(n481) );
  NAND2X0 U538 ( .IN1(n494), .IN2(n496), .QN(n495) );
  XNOR2X1 U539 ( .IN1(n497), .IN2(G2), .Q(n494) );
  AO21X1 U540 ( .IN1(G10), .IN2(n360), .IN3(n498), .Q(n496) );
  XOR2X1 U541 ( .IN1(keyinput8), .IN2(n499), .Q(n498) );
  NOR2X0 U542 ( .IN1(G10), .IN2(n360), .QN(n499) );
  INVX0 U543 ( .INP(G14), .ZN(n360) );
  INVX0 U544 ( .INP(n320), .ZN(n423) );
  XNOR3X1 U545 ( .IN1(n500), .IN2(n501), .IN3(n502), .Q(n320) );
  XNOR3X1 U546 ( .IN1(keyinput21), .IN2(G32), .IN3(G28), .Q(n502) );
  OA21X1 U547 ( .IN1(n503), .IN2(n504), .IN3(n505), .Q(n501) );
  XOR2X1 U548 ( .IN1(n506), .IN2(keyinput28), .Q(n505) );
  NAND2X0 U549 ( .IN1(n503), .IN2(n504), .QN(n506) );
  XOR2X1 U550 ( .IN1(n507), .IN2(n508), .Q(n504) );
  XOR2X1 U551 ( .IN1(n509), .IN2(keyinput2), .Q(n503) );
  NAND2X0 U552 ( .IN1(G40), .IN2(G41), .QN(n509) );
  OA21X1 U553 ( .IN1(G20), .IN2(G24), .IN3(n510), .Q(n500) );
  XOR2X1 U554 ( .IN1(n511), .IN2(keyinput4), .Q(n510) );
  NAND2X0 U555 ( .IN1(G24), .IN2(G20), .QN(n511) );
  NOR2X0 U556 ( .IN1(n305), .IN2(n408), .QN(n427) );
  INVX0 U557 ( .INP(n313), .ZN(n408) );
  AO21X1 U558 ( .IN1(n512), .IN2(n513), .IN3(n514), .Q(n313) );
  XOR2X1 U559 ( .IN1(n515), .IN2(keyinput32), .Q(n514) );
  NAND2X0 U560 ( .IN1(n516), .IN2(n513), .QN(n515) );
  NAND2X0 U561 ( .IN1(n516), .IN2(n512), .QN(n513) );
  AOI21X1 U562 ( .IN1(n517), .IN2(n518), .IN3(n519), .QN(n516) );
  XOR2X1 U563 ( .IN1(keyinput27), .IN2(n520), .Q(n519) );
  NOR2X0 U564 ( .IN1(n517), .IN2(n518), .QN(n520) );
  NAND2X0 U565 ( .IN1(G39), .IN2(G41), .QN(n518) );
  XNOR3X1 U566 ( .IN1(keyinput24), .IN2(n521), .IN3(n522), .Q(n517) );
  XNOR3X1 U567 ( .IN1(G23), .IN2(G19), .IN3(n523), .Q(n512) );
  XNOR2X1 U568 ( .IN1(G31), .IN2(G27), .Q(n523) );
  XNOR2X1 U569 ( .IN1(n524), .IN2(n525), .Q(n305) );
  XOR3X1 U570 ( .IN1(keyinput23), .IN2(keyinput19), .IN3(n526), .Q(n525) );
  XOR2X1 U571 ( .IN1(keyinput1), .IN2(n527), .Q(n526) );
  OA21X1 U572 ( .IN1(n528), .IN2(n529), .IN3(n530), .Q(n527) );
  XOR2X1 U573 ( .IN1(n531), .IN2(keyinput17), .Q(n530) );
  NAND3X0 U574 ( .IN1(n529), .IN2(n532), .IN3(n533), .QN(n531) );
  NAND2X0 U575 ( .IN1(G29), .IN2(n309), .QN(n532) );
  INVX0 U576 ( .INP(G25), .ZN(n309) );
  XNOR2X1 U577 ( .IN1(n334), .IN2(G17), .Q(n529) );
  INVX0 U578 ( .INP(G21), .ZN(n334) );
  OA21X1 U579 ( .IN1(G25), .IN2(n315), .IN3(n533), .Q(n528) );
  XOR2X1 U580 ( .IN1(n534), .IN2(keyinput11), .Q(n533) );
  NAND2X0 U581 ( .IN1(G25), .IN2(n315), .QN(n534) );
  INVX0 U582 ( .INP(G29), .ZN(n315) );
  XNOR3X1 U583 ( .IN1(n535), .IN2(n522), .IN3(n507), .Q(n524) );
  XOR2X1 U584 ( .IN1(n536), .IN2(n537), .Q(n507) );
  OA21X1 U585 ( .IN1(G5), .IN2(n497), .IN3(n538), .Q(n537) );
  XOR2X1 U586 ( .IN1(n539), .IN2(keyinput5), .Q(n538) );
  NAND2X0 U587 ( .IN1(G5), .IN2(n497), .QN(n539) );
  INVX0 U588 ( .INP(G6), .ZN(n497) );
  OA21X1 U589 ( .IN1(G7), .IN2(n540), .IN3(n541), .Q(n536) );
  XOR2X1 U590 ( .IN1(keyinput6), .IN2(n542), .Q(n541) );
  NOR2X0 U591 ( .IN1(G8), .IN2(n543), .QN(n542) );
  INVX0 U592 ( .INP(G7), .ZN(n543) );
  INVX0 U593 ( .INP(G8), .ZN(n540) );
  OAI21X1 U594 ( .IN1(n544), .IN2(n545), .IN3(n546), .QN(n522) );
  XNOR2X1 U595 ( .IN1(n547), .IN2(keyinput14), .Q(n546) );
  NAND2X0 U596 ( .IN1(n545), .IN2(n544), .QN(n547) );
  XNOR2X1 U597 ( .IN1(G1), .IN2(n394), .Q(n545) );
  INVX0 U598 ( .INP(G2), .ZN(n394) );
  XOR2X1 U599 ( .IN1(G4), .IN2(G3), .Q(n544) );
  NAND2X0 U600 ( .IN1(G37), .IN2(G41), .QN(n535) );
  XNOR2X1 U601 ( .IN1(n331), .IN2(keyinput34), .Q(n438) );
  INVX0 U602 ( .INP(n324), .ZN(n331) );
  MUX21X1 U603 ( .IN1(n548), .IN2(n549), .S(n550), .Q(n324) );
  XNOR3X1 U604 ( .IN1(keyinput20), .IN2(n416), .IN3(n551), .Q(n550) );
  XOR2X1 U605 ( .IN1(G26), .IN2(n552), .Q(n551) );
  OA21X1 U606 ( .IN1(G18), .IN2(n553), .IN3(n554), .Q(n552) );
  XOR2X1 U607 ( .IN1(n555), .IN2(keyinput12), .Q(n554) );
  NAND2X0 U608 ( .IN1(G18), .IN2(n553), .QN(n555) );
  INVX0 U609 ( .INP(G22), .ZN(n553) );
  INVX0 U610 ( .INP(G30), .ZN(n416) );
  NAND2X0 U611 ( .IN1(n556), .IN2(n557), .QN(n549) );
  AND2X1 U612 ( .IN1(n557), .IN2(n556), .Q(n548) );
  NAND3X0 U613 ( .IN1(G38), .IN2(G41), .IN3(n558), .QN(n556) );
  AO21X1 U614 ( .IN1(G38), .IN2(G41), .IN3(n558), .Q(n557) );
  XNOR2X1 U615 ( .IN1(n521), .IN2(n508), .Q(n558) );
  XNOR3X1 U616 ( .IN1(G14), .IN2(G13), .IN3(n559), .Q(n508) );
  XNOR2X1 U617 ( .IN1(G15), .IN2(G16), .Q(n559) );
  AOI21X1 U618 ( .IN1(n560), .IN2(n561), .IN3(n562), .QN(n521) );
  XOR2X1 U619 ( .IN1(keyinput15), .IN2(n563), .Q(n562) );
  NOR2X0 U620 ( .IN1(n560), .IN2(n561), .QN(n563) );
  XNOR2X1 U621 ( .IN1(n377), .IN2(G9), .Q(n561) );
  INVX0 U622 ( .INP(G10), .ZN(n377) );
  XNOR2X1 U623 ( .IN1(G12), .IN2(G11), .Q(n560) );
endmodule

