
module c7552 ( N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, 
        N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, 
        N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, 
        N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, 
        N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, 
        N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, 
        N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, 
        N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, 
        N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, 
        N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, 
        N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, 
        N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, 
        N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, 
        N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, 
        N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, 
        N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, 
        N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, 
        N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, 
        N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, 
        N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, 
        N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, 
        N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, 
        N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, 
        N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, 
        N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, 
        N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, 
        N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, 
        N11333, N11334, N11340, N11342, N241_O, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47,
         N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110,
         N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133,
         N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245,
         N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280,
         N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316,
         N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349,
         N352, N355, N358, N361, N364, N367, N382, N241_I, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507,
         N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543,
         N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567,
         N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884,
         N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490,
         N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111,
         N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576,
         N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713,
         N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760,
         N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840,
         N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908,
         N11333, N11334, N11340, N11342, N241_O;
  wire   N1, N106, N248, N251, N254, N257, N260, N263, N267, N274, N277, N280,
         N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316,
         N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349,
         N352, N355, N358, N361, N364, N241_I, N10102, N10706, N10759, N10837,
         N10839, N582, N1113, N1112, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089;
  assign N1490 = N1;
  assign N889 = N1;
  assign N388 = N1;
  assign N387 = N1;
  assign N945 = N106;
  assign N478 = N248;
  assign N643 = N251;
  assign N482 = N254;
  assign N484 = N257;
  assign N486 = N260;
  assign N489 = N263;
  assign N492 = N267;
  assign N501 = N274;
  assign N707 = N277;
  assign N505 = N280;
  assign N507 = N283;
  assign N509 = N286;
  assign N511 = N289;
  assign N513 = N293;
  assign N515 = N296;
  assign N517 = N299;
  assign N519 = N303;
  assign N535 = N307;
  assign N537 = N310;
  assign N539 = N313;
  assign N541 = N316;
  assign N543 = N319;
  assign N545 = N322;
  assign N547 = N325;
  assign N549 = N328;
  assign N551 = N331;
  assign N553 = N334;
  assign N556 = N337;
  assign N813 = N340;
  assign N559 = N343;
  assign N561 = N346;
  assign N563 = N349;
  assign N565 = N352;
  assign N567 = N355;
  assign N569 = N358;
  assign N571 = N361;
  assign N573 = N364;
  assign N241_O = N241_I;
  assign N10103 = N10102;
  assign N10104 = N10706;
  assign N10101 = N10759;
  assign N10838 = N10837;
  assign N10840 = N10839;
  assign N1114 = N582;
  assign N1111 = N582;
  assign N1489 = N1113;
  assign N1110 = N1112;

  INVX0 U1145 ( .INP(N18), .ZN(n1119) );
  INVX0 U1146 ( .INP(N18), .ZN(n1120) );
  INVX0 U1147 ( .INP(N18), .ZN(n1121) );
  INVX0 U1148 ( .INP(N18), .ZN(n1122) );
  OR2X1 U1149 ( .IN1(N5), .IN2(N57), .Q(N881) );
  INVX0 U1150 ( .INP(N15), .ZN(N582) );
  AND2X1 U1151 ( .IN1(N163), .IN2(N1), .Q(N1781) );
  XOR2X1 U1152 ( .IN1(n1123), .IN2(n1124), .Q(N11342) );
  NOR2X0 U1153 ( .IN1(keyinput125), .IN2(n1125), .QN(n1124) );
  MUX21X1 U1154 ( .IN1(n1126), .IN2(n1127), .S(n1128), .Q(n1125) );
  XOR2X1 U1155 ( .IN1(n1129), .IN2(n1130), .Q(n1127) );
  XNOR3X1 U1156 ( .IN1(keyinput123), .IN2(n1131), .IN3(n1132), .Q(n1130) );
  NOR2X0 U1157 ( .IN1(keyinput102), .IN2(n1133), .QN(n1132) );
  OA21X1 U1158 ( .IN1(n1134), .IN2(n1135), .IN3(n1136), .Q(n1133) );
  XOR2X1 U1159 ( .IN1(keyinput113), .IN2(n1137), .Q(n1136) );
  AND2X1 U1160 ( .IN1(n1134), .IN2(n1135), .Q(n1137) );
  XOR3X1 U1161 ( .IN1(n1138), .IN2(n1139), .IN3(n1140), .Q(n1135) );
  XNOR3X1 U1162 ( .IN1(n1141), .IN2(n1142), .IN3(n1143), .Q(n1129) );
  XOR3X1 U1163 ( .IN1(n1143), .IN2(n1144), .IN3(n1145), .Q(n1126) );
  MUX21X1 U1164 ( .IN1(n1146), .IN2(n1147), .S(n1148), .Q(n1145) );
  OA21X1 U1165 ( .IN1(n1142), .IN2(n1149), .IN3(n1134), .Q(n1148) );
  XNOR2X1 U1166 ( .IN1(keyinput114), .IN2(n1147), .Q(n1146) );
  XOR2X1 U1167 ( .IN1(n1150), .IN2(n1151), .Q(n1147) );
  NOR2X0 U1168 ( .IN1(keyinput104), .IN2(n1152), .QN(n1151) );
  XNOR2X1 U1169 ( .IN1(n1153), .IN2(n1154), .Q(n1152) );
  AO21X1 U1170 ( .IN1(n1140), .IN2(n1149), .IN3(keyinput73), .Q(n1153) );
  NAND2X0 U1171 ( .IN1(n1139), .IN2(n1155), .QN(n1150) );
  XNOR3X1 U1172 ( .IN1(n1156), .IN2(n1131), .IN3(n1157), .Q(n1144) );
  XNOR2X1 U1173 ( .IN1(n1158), .IN2(n1159), .Q(n1143) );
  OA21X1 U1174 ( .IN1(n1160), .IN2(n1161), .IN3(n1162), .Q(n1123) );
  MUX21X1 U1175 ( .IN1(n1163), .IN2(n1164), .S(n1165), .Q(n1162) );
  NAND2X0 U1176 ( .IN1(n1166), .IN2(n1161), .QN(n1164) );
  NAND2X0 U1177 ( .IN1(n1167), .IN2(n1168), .QN(n1163) );
  XNOR2X1 U1178 ( .IN1(keyinput90), .IN2(n1161), .Q(n1168) );
  MUX21X1 U1179 ( .IN1(n1167), .IN2(n1166), .S(n1165), .Q(n1160) );
  XNOR3X1 U1180 ( .IN1(n1169), .IN2(n1170), .IN3(n1171), .Q(n1166) );
  XNOR2X1 U1181 ( .IN1(n1172), .IN2(n1173), .Q(n1171) );
  AOI21X1 U1182 ( .IN1(n1174), .IN2(n1175), .IN3(n1176), .QN(n1173) );
  MUX21X1 U1183 ( .IN1(n1177), .IN2(n1178), .S(n1179), .Q(n1170) );
  NOR2X0 U1184 ( .IN1(n1175), .IN2(n1178), .QN(n1177) );
  XOR2X1 U1185 ( .IN1(n1180), .IN2(n1181), .Q(n1167) );
  XNOR2X1 U1186 ( .IN1(n1182), .IN2(n1169), .Q(n1181) );
  XNOR2X1 U1187 ( .IN1(n1183), .IN2(n1184), .Q(n1169) );
  XNOR3X1 U1188 ( .IN1(n1178), .IN2(n1172), .IN3(n1176), .Q(n1180) );
  OA21X1 U1189 ( .IN1(n1185), .IN2(n1186), .IN3(n1187), .Q(N11340) );
  XOR2X1 U1190 ( .IN1(n1188), .IN2(keyinput127), .Q(n1187) );
  NAND2X0 U1191 ( .IN1(n1189), .IN2(n1186), .QN(n1188) );
  XNOR2X1 U1192 ( .IN1(n1185), .IN2(keyinput126), .Q(n1189) );
  AO22X1 U1193 ( .IN1(n1190), .IN2(n1191), .IN3(n1192), .IN4(n1193), .Q(n1186)
         );
  XOR2X1 U1194 ( .IN1(n1194), .IN2(n1195), .Q(n1192) );
  XNOR3X1 U1195 ( .IN1(n1196), .IN2(n1197), .IN3(n1198), .Q(n1195) );
  XNOR3X1 U1196 ( .IN1(n1199), .IN2(n1200), .IN3(n1201), .Q(n1194) );
  MUX21X1 U1197 ( .IN1(n1202), .IN2(n1203), .S(n1204), .Q(n1201) );
  AO21X1 U1198 ( .IN1(n1205), .IN2(n1206), .IN3(n1207), .Q(n1203) );
  OA21X1 U1199 ( .IN1(n1208), .IN2(n1209), .IN3(n1210), .Q(n1202) );
  NAND2X0 U1200 ( .IN1(keyinput108), .IN2(n1211), .QN(n1200) );
  XNOR3X1 U1201 ( .IN1(n1212), .IN2(n1197), .IN3(n1199), .Q(n1191) );
  XOR3X1 U1202 ( .IN1(n1209), .IN2(n1213), .IN3(n1214), .Q(n1199) );
  OA21X1 U1203 ( .IN1(n1196), .IN2(n1215), .IN3(n1216), .Q(n1212) );
  XOR2X1 U1204 ( .IN1(n1217), .IN2(keyinput118), .Q(n1216) );
  NAND2X0 U1205 ( .IN1(n1215), .IN2(n1196), .QN(n1217) );
  XNOR3X1 U1206 ( .IN1(n1218), .IN2(n1219), .IN3(n1220), .Q(n1215) );
  NAND2X0 U1207 ( .IN1(keyinput106), .IN2(n1221), .QN(n1220) );
  XOR3X1 U1208 ( .IN1(keyinput105), .IN2(n1222), .IN3(n1223), .Q(n1221) );
  OA21X1 U1209 ( .IN1(n1219), .IN2(n1209), .IN3(n1210), .Q(n1223) );
  OA21X1 U1210 ( .IN1(n1196), .IN2(n1197), .IN3(n1211), .Q(n1219) );
  INVX0 U1211 ( .INP(n1224), .ZN(n1197) );
  NOR2X0 U1212 ( .IN1(n1225), .IN2(n1198), .QN(n1218) );
  NAND4X0 U1213 ( .IN1(n1226), .IN2(n1227), .IN3(n1228), .IN4(n1229), .QN(
        n1198) );
  NAND2X0 U1214 ( .IN1(n1230), .IN2(n1204), .QN(n1226) );
  XOR2X1 U1215 ( .IN1(keyinput124), .IN2(n1231), .Q(n1185) );
  OA22X1 U1216 ( .IN1(n1232), .IN2(n1233), .IN3(n1234), .IN4(n1235), .Q(n1231)
         );
  XOR3X1 U1217 ( .IN1(n1236), .IN2(n1237), .IN3(n1238), .Q(n1235) );
  XNOR2X1 U1218 ( .IN1(n1239), .IN2(n1240), .Q(n1238) );
  NAND3X0 U1219 ( .IN1(n1241), .IN2(n1242), .IN3(n1243), .QN(n1239) );
  XOR2X1 U1220 ( .IN1(n1244), .IN2(keyinput78), .Q(n1243) );
  OR2X1 U1221 ( .IN1(n1245), .IN2(n1246), .Q(n1244) );
  OR2X1 U1222 ( .IN1(n1247), .IN2(n1246), .Q(n1241) );
  XNOR3X1 U1223 ( .IN1(n1248), .IN2(n1249), .IN3(n1250), .Q(n1236) );
  XNOR2X1 U1224 ( .IN1(n1251), .IN2(n1252), .Q(n1250) );
  OA22X1 U1225 ( .IN1(n1253), .IN2(n1254), .IN3(n1255), .IN4(n1256), .Q(n1234)
         );
  INVX0 U1226 ( .INP(n1193), .ZN(n1255) );
  OA21X1 U1227 ( .IN1(n1257), .IN2(n1246), .IN3(n1258), .Q(n1233) );
  XOR2X1 U1228 ( .IN1(n1259), .IN2(keyinput122), .Q(n1258) );
  NAND2X0 U1229 ( .IN1(n1257), .IN2(n1246), .QN(n1259) );
  XOR3X1 U1230 ( .IN1(n1260), .IN2(n1261), .IN3(n1262), .Q(n1257) );
  XOR2X1 U1231 ( .IN1(n1237), .IN2(n1263), .Q(n1262) );
  OA21X1 U1232 ( .IN1(n1246), .IN2(n1264), .IN3(n1265), .Q(n1263) );
  INVX0 U1233 ( .INP(n1252), .ZN(n1246) );
  XOR3X1 U1234 ( .IN1(keyinput87), .IN2(n1248), .IN3(n1249), .Q(n1261) );
  MUX21X1 U1235 ( .IN1(n1240), .IN2(n1266), .S(n1267), .Q(n1260) );
  NOR2X0 U1236 ( .IN1(n1268), .IN2(n1240), .QN(n1266) );
  AOI22X1 U1237 ( .IN1(n1254), .IN2(n1190), .IN3(n1256), .IN4(n1193), .QN(
        n1232) );
  XOR2X1 U1238 ( .IN1(n1253), .IN2(keyinput112), .Q(n1193) );
  INVX0 U1239 ( .INP(n1190), .ZN(n1253) );
  MUX21X1 U1240 ( .IN1(n1269), .IN2(n1270), .S(keyinput109), .Q(n1190) );
  OAI21X1 U1241 ( .IN1(n1271), .IN2(n1272), .IN3(n1165), .QN(n1270) );
  AO21X1 U1242 ( .IN1(n1225), .IN2(n1273), .IN3(n1256), .Q(n1254) );
  INVX0 U1243 ( .INP(n1274), .ZN(n1256) );
  XOR2X1 U1244 ( .IN1(n1275), .IN2(n1276), .Q(N11334) );
  MUX21X1 U1245 ( .IN1(n1277), .IN2(n1278), .S(n1279), .Q(n1276) );
  XOR3X1 U1246 ( .IN1(n1280), .IN2(n1281), .IN3(n1282), .Q(n1278) );
  XNOR3X1 U1247 ( .IN1(n1283), .IN2(n1284), .IN3(n1285), .Q(n1282) );
  MUX21X1 U1248 ( .IN1(n1286), .IN2(n1287), .S(n1288), .Q(n1285) );
  AOI21X1 U1249 ( .IN1(n1289), .IN2(n1290), .IN3(n1287), .QN(n1286) );
  AO21X1 U1250 ( .IN1(n1291), .IN2(n1289), .IN3(n1292), .Q(n1287) );
  XOR2X1 U1251 ( .IN1(n1293), .IN2(n1294), .Q(n1281) );
  XNOR2X1 U1252 ( .IN1(n1295), .IN2(n1296), .Q(n1280) );
  XOR2X1 U1253 ( .IN1(n1297), .IN2(n1298), .Q(n1277) );
  XOR3X1 U1254 ( .IN1(n1283), .IN2(n1284), .IN3(n1299), .Q(n1298) );
  XOR2X1 U1255 ( .IN1(n1300), .IN2(n1301), .Q(n1299) );
  NOR2X0 U1256 ( .IN1(n1302), .IN2(n1303), .QN(n1301) );
  AOI21X1 U1257 ( .IN1(n1289), .IN2(n1304), .IN3(n1292), .QN(n1300) );
  XOR2X1 U1258 ( .IN1(n1289), .IN2(n1305), .Q(n1284) );
  XNOR3X1 U1259 ( .IN1(n1306), .IN2(n1290), .IN3(n1307), .Q(n1297) );
  XNOR2X1 U1260 ( .IN1(n1308), .IN2(n1304), .Q(n1307) );
  OA21X1 U1261 ( .IN1(n1309), .IN2(n1310), .IN3(n1293), .Q(n1308) );
  OA21X1 U1262 ( .IN1(n1309), .IN2(n1294), .IN3(n1311), .Q(n1293) );
  MUX21X1 U1263 ( .IN1(n1312), .IN2(n1313), .S(n1314), .Q(n1275) );
  XNOR2X1 U1264 ( .IN1(n1315), .IN2(n1316), .Q(n1313) );
  XNOR2X1 U1265 ( .IN1(n1315), .IN2(n1317), .Q(n1312) );
  AO21X1 U1266 ( .IN1(n1318), .IN2(n1319), .IN3(n1320), .Q(n1315) );
  XNOR3X1 U1267 ( .IN1(n1321), .IN2(n1322), .IN3(n1323), .Q(N11333) );
  MUX21X1 U1268 ( .IN1(n1324), .IN2(n1325), .S(n1326), .Q(n1322) );
  XNOR3X1 U1269 ( .IN1(n1327), .IN2(n1328), .IN3(n1329), .Q(n1325) );
  NOR2X0 U1270 ( .IN1(keyinput81), .IN2(n1330), .QN(n1327) );
  XOR3X1 U1271 ( .IN1(n1331), .IN2(n1332), .IN3(n1333), .Q(n1330) );
  NAND2X0 U1272 ( .IN1(n1334), .IN2(n1335), .QN(n1333) );
  XOR2X1 U1273 ( .IN1(keyinput68), .IN2(n1336), .Q(n1335) );
  XOR2X1 U1274 ( .IN1(n1337), .IN2(n1338), .Q(n1332) );
  NOR2X0 U1275 ( .IN1(keyinput98), .IN2(n1339), .QN(n1337) );
  NOR2X0 U1276 ( .IN1(n1340), .IN2(n1341), .QN(n1331) );
  XNOR3X1 U1277 ( .IN1(keyinput120), .IN2(n1342), .IN3(n1343), .Q(n1324) );
  OA21X1 U1278 ( .IN1(n1344), .IN2(n1345), .IN3(n1346), .Q(n1342) );
  XOR2X1 U1279 ( .IN1(keyinput117), .IN2(n1347), .Q(n1346) );
  AND2X1 U1280 ( .IN1(n1344), .IN2(n1345), .Q(n1347) );
  XNOR3X1 U1281 ( .IN1(n1348), .IN2(n1341), .IN3(n1349), .Q(n1345) );
  XNOR2X1 U1282 ( .IN1(n1334), .IN2(n1338), .Q(n1349) );
  OA21X1 U1283 ( .IN1(n1343), .IN2(n1350), .IN3(n1351), .Q(n1334) );
  INVX0 U1284 ( .INP(n1328), .ZN(n1343) );
  OA21X1 U1285 ( .IN1(n1352), .IN2(n1353), .IN3(n1354), .Q(n1321) );
  MUX21X1 U1286 ( .IN1(n1355), .IN2(n1356), .S(n1357), .Q(n1354) );
  NAND2X0 U1287 ( .IN1(n1358), .IN2(n1352), .QN(n1356) );
  XNOR2X1 U1288 ( .IN1(n1357), .IN2(n1358), .Q(n1353) );
  XOR2X1 U1289 ( .IN1(n1359), .IN2(n1360), .Q(n1357) );
  MUX21X1 U1290 ( .IN1(n1361), .IN2(n1362), .S(n1363), .Q(n1360) );
  XOR3X1 U1291 ( .IN1(n1364), .IN2(n1365), .IN3(n1366), .Q(n1362) );
  XNOR2X1 U1292 ( .IN1(n1367), .IN2(n1368), .Q(n1366) );
  NOR2X0 U1293 ( .IN1(keyinput121), .IN2(n1369), .QN(n1368) );
  OA21X1 U1294 ( .IN1(n1355), .IN2(n1370), .IN3(n1371), .Q(n1365) );
  OA21X1 U1295 ( .IN1(n1372), .IN2(n1373), .IN3(n1374), .Q(n1364) );
  XOR2X1 U1296 ( .IN1(n1375), .IN2(keyinput103), .Q(n1374) );
  NAND3X0 U1297 ( .IN1(n1376), .IN2(n1370), .IN3(n1373), .QN(n1375) );
  XOR2X1 U1298 ( .IN1(n1377), .IN2(n1378), .Q(n1373) );
  NOR2X0 U1299 ( .IN1(n1379), .IN2(n1380), .QN(n1378) );
  OA21X1 U1300 ( .IN1(n1381), .IN2(n1382), .IN3(n1383), .Q(n1380) );
  NAND2X0 U1301 ( .IN1(N277), .IN2(n1384), .QN(n1377) );
  NOR2X0 U1302 ( .IN1(n1381), .IN2(n1382), .QN(n1372) );
  NOR2X0 U1303 ( .IN1(keyinput82), .IN2(n1385), .QN(n1361) );
  XNOR3X1 U1304 ( .IN1(n1386), .IN2(n1376), .IN3(n1387), .Q(n1385) );
  XNOR3X1 U1305 ( .IN1(n1369), .IN2(n1371), .IN3(n1388), .Q(n1387) );
  OA21X1 U1306 ( .IN1(n1358), .IN2(n1389), .IN3(n1390), .Q(n1388) );
  XNOR2X1 U1307 ( .IN1(n1391), .IN2(n1392), .Q(n1390) );
  OA21X1 U1308 ( .IN1(n1358), .IN2(n1393), .IN3(n1394), .Q(n1392) );
  INVX0 U1309 ( .INP(n1383), .ZN(n1358) );
  NAND3X0 U1310 ( .IN1(N134), .IN2(N133), .IN3(n1395), .QN(N1113) );
  XNOR2X1 U1311 ( .IN1(N5), .IN2(keyinput0), .Q(n1395) );
  NAND2X0 U1312 ( .IN1(N242), .IN2(n1396), .QN(N1112) );
  INVX0 U1313 ( .INP(N5), .ZN(n1396) );
  XNOR2X1 U1314 ( .IN1(n1249), .IN2(n1397), .Q(N10908) );
  XOR2X1 U1315 ( .IN1(n1248), .IN2(n1398), .Q(N10907) );
  OA21X1 U1316 ( .IN1(n1251), .IN2(n1399), .IN3(n1267), .Q(n1398) );
  MUX21X1 U1317 ( .IN1(n1400), .IN2(n1401), .S(n1399), .Q(N10906) );
  XOR2X1 U1318 ( .IN1(n1402), .IN2(n1403), .Q(n1401) );
  XOR2X1 U1319 ( .IN1(n1404), .IN2(n1403), .Q(n1400) );
  NAND2X0 U1320 ( .IN1(n1405), .IN2(n1406), .QN(N10905) );
  OR3X1 U1321 ( .IN1(n1399), .IN2(n1407), .IN3(n1408), .Q(n1406) );
  MUX21X1 U1322 ( .IN1(n1409), .IN2(n1410), .S(n1237), .Q(n1405) );
  NAND2X0 U1323 ( .IN1(n1411), .IN2(n1242), .QN(n1410) );
  AO22X1 U1324 ( .IN1(n1411), .IN2(n1242), .IN3(n1407), .IN4(n1397), .Q(n1409)
         );
  INVX0 U1325 ( .INP(n1399), .ZN(n1397) );
  AO21X1 U1326 ( .IN1(n1412), .IN2(n1413), .IN3(n1414), .Q(n1399) );
  NOR2X0 U1327 ( .IN1(n1408), .IN2(n1237), .QN(n1407) );
  NAND2X0 U1328 ( .IN1(n1403), .IN2(n1402), .QN(n1411) );
  OR2X1 U1329 ( .IN1(n1404), .IN2(n1268), .Q(n1402) );
  XNOR2X1 U1330 ( .IN1(n1224), .IN2(n1415), .Q(N10871) );
  XNOR2X1 U1331 ( .IN1(n1205), .IN2(n1416), .Q(N10870) );
  XOR3X1 U1332 ( .IN1(keyinput119), .IN2(n1417), .IN3(n1418), .Q(N10869) );
  NAND2X0 U1333 ( .IN1(keyinput116), .IN2(n1419), .QN(n1418) );
  OA21X1 U1334 ( .IN1(n1209), .IN2(n1416), .IN3(n1210), .Q(n1417) );
  AO21X1 U1335 ( .IN1(n1415), .IN2(n1208), .IN3(n1420), .Q(n1416) );
  OA21X1 U1336 ( .IN1(n1196), .IN2(n1421), .IN3(n1422), .Q(n1415) );
  INVX0 U1337 ( .INP(n1423), .ZN(n1196) );
  XOR2X1 U1338 ( .IN1(n1413), .IN2(n1412), .Q(N10868) );
  AO21X1 U1339 ( .IN1(n1225), .IN2(n1424), .IN3(n1425), .Q(n1413) );
  XNOR2X1 U1340 ( .IN1(n1423), .IN2(n1421), .Q(N10827) );
  INVX0 U1341 ( .INP(n1424), .ZN(n1421) );
  NAND3X0 U1342 ( .IN1(n1426), .IN2(n1427), .IN3(n1428), .QN(n1424) );
  NAND2X0 U1343 ( .IN1(n1429), .IN2(n1430), .QN(n1428) );
  XOR2X1 U1344 ( .IN1(keyinput89), .IN2(n1272), .Q(n1429) );
  XNOR2X1 U1345 ( .IN1(n1431), .IN2(n1319), .Q(N10839) );
  XOR2X1 U1346 ( .IN1(n1432), .IN2(n1318), .Q(N10837) );
  AOI21X1 U1347 ( .IN1(n1316), .IN2(n1431), .IN3(n1433), .QN(n1432) );
  XNOR2X1 U1348 ( .IN1(n1434), .IN2(n1435), .Q(N10763) );
  AO21X1 U1349 ( .IN1(n1436), .IN2(n1437), .IN3(n1438), .Q(N10762) );
  XOR2X1 U1350 ( .IN1(n1439), .IN2(keyinput115), .Q(n1438) );
  NAND3X0 U1351 ( .IN1(n1440), .IN2(n1441), .IN3(n1434), .QN(n1439) );
  OR2X1 U1352 ( .IN1(n1442), .IN2(n1443), .Q(n1440) );
  XOR3X1 U1353 ( .IN1(keyinput93), .IN2(n1339), .IN3(n1442), .Q(n1436) );
  XNOR2X1 U1354 ( .IN1(n1444), .IN2(n1445), .Q(N10761) );
  NAND3X0 U1355 ( .IN1(n1441), .IN2(n1446), .IN3(n1447), .QN(n1444) );
  NAND2X0 U1356 ( .IN1(n1437), .IN2(n1448), .QN(n1447) );
  MUX21X1 U1357 ( .IN1(n1449), .IN2(n1450), .S(n1437), .Q(N10760) );
  XNOR3X1 U1358 ( .IN1(keyinput75), .IN2(n1451), .IN3(n1452), .Q(n1450) );
  AOI21X1 U1359 ( .IN1(n1448), .IN2(n1453), .IN3(n1454), .QN(n1451) );
  NAND3X0 U1360 ( .IN1(n1455), .IN2(n1446), .IN3(n1441), .QN(n1448) );
  OA21X1 U1361 ( .IN1(n1323), .IN2(n1456), .IN3(n1457), .Q(n1449) );
  NAND4X0 U1362 ( .IN1(n1458), .IN2(n1459), .IN3(n1460), .IN4(n1461), .QN(
        N10729) );
  NOR3X0 U1363 ( .IN1(N10576), .IN2(N883), .IN3(N882), .QN(n1461) );
  NAND4X0 U1364 ( .IN1(N240), .IN2(N228), .IN3(N184), .IN4(N150), .QN(N882) );
  NAND4X0 U1365 ( .IN1(N230), .IN2(N218), .IN3(N210), .IN4(N152), .QN(N883) );
  XOR2X1 U1366 ( .IN1(keyinput6), .IN2(n1462), .Q(n1460) );
  NOR2X0 U1367 ( .IN1(N885), .IN2(N884), .QN(n1462) );
  NAND4X0 U1368 ( .IN1(N186), .IN2(N185), .IN3(N183), .IN4(N182), .QN(N884) );
  NAND4X0 U1369 ( .IN1(N199), .IN2(N188), .IN3(N172), .IN4(N162), .QN(N885) );
  INVX0 U1370 ( .INP(N10575), .ZN(n1459) );
  INVX0 U1371 ( .INP(N10574), .ZN(n1458) );
  XNOR2X1 U1372 ( .IN1(n1463), .IN2(n1296), .Q(N10718) );
  NAND2X0 U1373 ( .IN1(n1464), .IN2(n1288), .QN(n1463) );
  XOR2X1 U1374 ( .IN1(n1465), .IN2(keyinput110), .Q(n1464) );
  NAND2X0 U1375 ( .IN1(n1466), .IN2(n1467), .QN(n1465) );
  XOR2X1 U1376 ( .IN1(n1468), .IN2(n1469), .Q(N10717) );
  XNOR2X1 U1377 ( .IN1(n1470), .IN2(n1295), .Q(N10716) );
  XNOR2X1 U1378 ( .IN1(n1471), .IN2(n1472), .Q(N10715) );
  OA21X1 U1379 ( .IN1(n1470), .IN2(n1306), .IN3(n1473), .Q(n1472) );
  AOI21X1 U1380 ( .IN1(n1469), .IN2(n1468), .IN3(n1292), .QN(n1470) );
  INVX0 U1381 ( .INP(n1474), .ZN(n1292) );
  XNOR2X1 U1382 ( .IN1(n1475), .IN2(n1476), .Q(N10714) );
  XNOR2X1 U1383 ( .IN1(n1477), .IN2(n1478), .Q(N10713) );
  NOR2X0 U1384 ( .IN1(n1479), .IN2(n1382), .QN(n1478) );
  XOR2X1 U1385 ( .IN1(n1480), .IN2(n1352), .Q(N10712) );
  NAND3X0 U1386 ( .IN1(n1481), .IN2(n1394), .IN3(n1482), .QN(n1480) );
  XOR2X1 U1387 ( .IN1(n1483), .IN2(keyinput70), .Q(n1482) );
  OR2X1 U1388 ( .IN1(n1393), .IN2(n1484), .Q(n1483) );
  OR3X1 U1389 ( .IN1(n1476), .IN2(n1484), .IN3(n1369), .Q(n1481) );
  OA21X1 U1390 ( .IN1(n1386), .IN2(n1485), .IN3(n1486), .Q(n1476) );
  XNOR2X1 U1391 ( .IN1(n1359), .IN2(n1487), .Q(N10711) );
  OA21X1 U1392 ( .IN1(n1488), .IN2(n1489), .IN3(n1490), .Q(n1487) );
  OA21X1 U1393 ( .IN1(n1484), .IN2(n1491), .IN3(n1492), .Q(n1489) );
  INVX0 U1394 ( .INP(n1477), .ZN(n1484) );
  AND4X1 U1395 ( .IN1(n1477), .IN2(n1491), .IN3(n1352), .IN4(n1493), .Q(n1488)
         );
  NAND2X0 U1396 ( .IN1(n1352), .IN2(n1494), .QN(n1491) );
  NAND3X0 U1397 ( .IN1(n1393), .IN2(n1495), .IN3(n1496), .QN(n1494) );
  NAND2X0 U1398 ( .IN1(n1493), .IN2(n1492), .QN(n1496) );
  INVX0 U1399 ( .INP(keyinput69), .ZN(n1492) );
  AO21X1 U1400 ( .IN1(n1320), .IN2(n1314), .IN3(n1497), .Q(N10706) );
  AO21X1 U1401 ( .IN1(n1305), .IN2(n1498), .IN3(n1499), .Q(n1314) );
  NAND2X0 U1402 ( .IN1(n1311), .IN2(n1500), .QN(n1498) );
  NAND3X0 U1403 ( .IN1(n1501), .IN2(n1304), .IN3(n1502), .QN(n1500) );
  INVX0 U1404 ( .INP(n1309), .ZN(n1502) );
  NAND2X0 U1405 ( .IN1(n1295), .IN2(n1289), .QN(n1309) );
  AO21X1 U1406 ( .IN1(N106), .IN2(n1503), .IN3(n1504), .Q(n1289) );
  XOR2X1 U1407 ( .IN1(n1505), .IN2(keyinput46), .Q(n1504) );
  OR2X1 U1408 ( .IN1(n1503), .IN2(N106), .Q(n1505) );
  NAND2X0 U1409 ( .IN1(n1294), .IN2(n1310), .QN(n1304) );
  OR2X1 U1410 ( .IN1(n1283), .IN2(n1296), .Q(n1310) );
  XOR2X1 U1411 ( .IN1(n1506), .IN2(n1302), .Q(n1283) );
  NAND2X0 U1412 ( .IN1(keyinput10), .IN2(n1303), .QN(n1506) );
  NAND2X0 U1413 ( .IN1(n1279), .IN2(n1294), .QN(n1501) );
  AOI221X1 U1414 ( .IN1(keyinput67), .IN2(n1507), .IN3(n1323), .IN4(n1508), 
        .IN5(n1509), .QN(n1279) );
  AO222X1 U1415 ( .IN1(n1328), .IN2(n1341), .IN3(n1336), .IN4(n1326), .IN5(
        n1454), .IN6(n1510), .Q(n1508) );
  INVX0 U1416 ( .INP(keyinput67), .ZN(n1510) );
  AO21X1 U1417 ( .IN1(n1359), .IN2(n1511), .IN3(n1512), .Q(n1326) );
  NAND2X0 U1418 ( .IN1(n1371), .IN2(n1513), .QN(n1511) );
  NAND3X0 U1419 ( .IN1(n1514), .IN2(n1363), .IN3(n1381), .QN(n1513) );
  AO22X1 U1420 ( .IN1(n1515), .IN2(n1516), .IN3(n1237), .IN4(n1517), .Q(n1363)
         );
  NAND2X0 U1421 ( .IN1(n1265), .IN2(n1518), .QN(n1517) );
  NAND3X0 U1422 ( .IN1(n1252), .IN2(n1519), .IN3(n1268), .QN(n1518) );
  NAND2X0 U1423 ( .IN1(n1274), .IN2(n1520), .QN(n1519) );
  NAND3X0 U1424 ( .IN1(n1273), .IN2(n1269), .IN3(n1225), .QN(n1520) );
  AO21X1 U1425 ( .IN1(n1272), .IN2(n1165), .IN3(n1271), .Q(n1269) );
  AO21X1 U1426 ( .IN1(n1184), .IN2(n1176), .IN3(n1521), .Q(n1271) );
  XOR2X1 U1427 ( .IN1(n1427), .IN2(keyinput35), .Q(n1521) );
  AO21X1 U1428 ( .IN1(n1174), .IN2(n1178), .IN3(n1522), .Q(n1176) );
  AO21X1 U1429 ( .IN1(n1523), .IN2(n1182), .IN3(n1524), .Q(n1178) );
  AO221X1 U1430 ( .IN1(n1141), .IN2(n1525), .IN3(n1526), .IN4(n1157), .IN5(
        n1527), .Q(n1165) );
  INVX0 U1431 ( .INP(n1134), .ZN(n1525) );
  OA21X1 U1432 ( .IN1(n1142), .IN2(n1140), .IN3(n1528), .Q(n1134) );
  OA21X1 U1433 ( .IN1(n1529), .IN2(n1139), .IN3(n1530), .Q(n1140) );
  OA21X1 U1434 ( .IN1(n1138), .IN2(n1159), .IN3(n1531), .Q(n1139) );
  INVX0 U1435 ( .INP(n1532), .ZN(n1531) );
  INVX0 U1436 ( .INP(n1157), .ZN(n1142) );
  XOR2X1 U1437 ( .IN1(N319), .IN2(n1533), .Q(n1157) );
  INVX0 U1438 ( .INP(n1214), .ZN(n1273) );
  OA21X1 U1439 ( .IN1(n1534), .IN2(n1214), .IN3(n1535), .Q(n1274) );
  INVX0 U1440 ( .INP(n1414), .ZN(n1535) );
  XOR2X1 U1441 ( .IN1(N352), .IN2(n1536), .Q(n1214) );
  NOR2X0 U1442 ( .IN1(keyinput14), .IN2(n1537), .QN(n1536) );
  OA21X1 U1443 ( .IN1(n1538), .IN2(n1213), .IN3(n1229), .Q(n1534) );
  INVX0 U1444 ( .INP(n1419), .ZN(n1213) );
  OA21X1 U1445 ( .IN1(n1209), .IN2(n1211), .IN3(n1210), .Q(n1538) );
  OAI21X1 U1446 ( .IN1(n1204), .IN2(n1539), .IN3(n1206), .QN(n1211) );
  INVX0 U1447 ( .INP(n1420), .ZN(n1206) );
  NOR2X0 U1448 ( .IN1(n1224), .IN2(n1539), .QN(n1420) );
  XOR2X1 U1449 ( .IN1(n1422), .IN2(keyinput39), .Q(n1204) );
  INVX0 U1450 ( .INP(n1205), .ZN(n1209) );
  AOI21X1 U1451 ( .IN1(n1252), .IN2(n1240), .IN3(n1540), .QN(n1265) );
  NAND2X0 U1452 ( .IN1(n1245), .IN2(n1247), .QN(n1240) );
  INVX0 U1453 ( .INP(n1355), .ZN(n1514) );
  OA21X1 U1454 ( .IN1(n1355), .IN2(n1376), .IN3(n1490), .Q(n1371) );
  NAND2X0 U1455 ( .IN1(n1352), .IN2(n1383), .QN(n1355) );
  AO22X1 U1456 ( .IN1(n1541), .IN2(n1542), .IN3(n1543), .IN4(n1544), .Q(n1383)
         );
  NOR2X0 U1457 ( .IN1(keyinput13), .IN2(n1379), .QN(n1543) );
  OR2X1 U1458 ( .IN1(n1394), .IN2(keyinput13), .Q(n1542) );
  AND2X1 U1459 ( .IN1(n1340), .IN2(n1328), .Q(n1336) );
  AND2X1 U1460 ( .IN1(n1329), .IN2(n1338), .Q(n1340) );
  XOR2X1 U1461 ( .IN1(n1435), .IN2(keyinput55), .Q(n1338) );
  INVX0 U1462 ( .INP(n1344), .ZN(n1329) );
  INVX0 U1463 ( .INP(n1350), .ZN(n1341) );
  OA21X1 U1464 ( .IN1(n1348), .IN2(n1344), .IN3(n1446), .Q(n1350) );
  XOR2X1 U1465 ( .IN1(N296), .IN2(n1545), .Q(n1344) );
  NOR2X0 U1466 ( .IN1(n1546), .IN2(keyinput12), .QN(n1545) );
  AO22X1 U1467 ( .IN1(n1547), .IN2(n1548), .IN3(n1549), .IN4(n1351), .Q(n1328)
         );
  NOR2X0 U1468 ( .IN1(keyinput30), .IN2(N299), .QN(n1549) );
  OR2X1 U1469 ( .IN1(n1351), .IN2(keyinput30), .Q(n1547) );
  INVX0 U1470 ( .INP(n1454), .ZN(n1351) );
  NAND2X0 U1471 ( .IN1(n1323), .IN2(n1454), .QN(n1507) );
  NAND2X0 U1472 ( .IN1(n1550), .IN2(n1551), .QN(n1305) );
  XNOR2X1 U1473 ( .IN1(keyinput45), .IN2(n1552), .Q(n1551) );
  XOR2X1 U1474 ( .IN1(n1553), .IN2(keyinput27), .Q(n1550) );
  AO21X1 U1475 ( .IN1(n1554), .IN2(n1555), .IN3(n1556), .Q(N10704) );
  XOR2X1 U1476 ( .IN1(n1557), .IN2(n1558), .Q(n1556) );
  NOR2X0 U1477 ( .IN1(n1559), .IN2(keyinput95), .QN(n1558) );
  INVX0 U1478 ( .INP(n1555), .ZN(n1559) );
  NAND2X0 U1479 ( .IN1(n1560), .IN2(n1561), .QN(n1555) );
  NAND4X0 U1480 ( .IN1(n1562), .IN2(n1563), .IN3(n1564), .IN4(n1565), .QN(
        n1561) );
  NAND2X0 U1481 ( .IN1(n1566), .IN2(n1567), .QN(n1564) );
  AO21X1 U1482 ( .IN1(n1568), .IN2(n1569), .IN3(n1570), .Q(n1567) );
  XOR2X1 U1483 ( .IN1(n1466), .IN2(n1467), .Q(N10641) );
  XNOR2X1 U1484 ( .IN1(n1367), .IN2(n1485), .Q(N10632) );
  AO21X1 U1485 ( .IN1(n1571), .IN2(n1572), .IN3(n1573), .Q(N10628) );
  XNOR2X1 U1486 ( .IN1(n1574), .IN2(n1575), .Q(n1573) );
  NOR2X0 U1487 ( .IN1(n1576), .IN2(keyinput51), .QN(n1575) );
  INVX0 U1488 ( .INP(n1572), .ZN(n1576) );
  NAND2X0 U1489 ( .IN1(n1577), .IN2(n1578), .QN(n1572) );
  XNOR2X1 U1490 ( .IN1(n1579), .IN2(keyinput83), .Q(n1577) );
  INVX0 U1491 ( .INP(n1580), .ZN(n1571) );
  NAND4X0 U1492 ( .IN1(n1581), .IN2(n1582), .IN3(n1583), .IN4(n1584), .QN(
        N10576) );
  XNOR3X1 U1493 ( .IN1(n1585), .IN2(n1586), .IN3(n1587), .Q(n1584) );
  AO21X1 U1494 ( .IN1(N164), .IN2(n1588), .IN3(n1589), .Q(n1587) );
  OA21X1 U1495 ( .IN1(n1590), .IN2(n1591), .IN3(n1592), .Q(n1586) );
  XOR2X1 U1496 ( .IN1(keyinput88), .IN2(n1593), .Q(n1592) );
  NOR2X0 U1497 ( .IN1(n1594), .IN2(n1595), .QN(n1593) );
  XNOR2X1 U1498 ( .IN1(n1596), .IN2(n1597), .Q(n1595) );
  INVX0 U1499 ( .INP(n1594), .ZN(n1591) );
  XOR2X1 U1500 ( .IN1(n1598), .IN2(n1599), .Q(n1594) );
  XOR2X1 U1501 ( .IN1(n1597), .IN2(n1596), .Q(n1590) );
  NOR3X0 U1502 ( .IN1(N170), .IN2(n1600), .IN3(n1120), .QN(n1596) );
  AO21X1 U1503 ( .IN1(n1601), .IN2(n1602), .IN3(n1603), .Q(n1597) );
  XOR2X1 U1504 ( .IN1(keyinput47), .IN2(n1604), .Q(n1603) );
  NOR2X0 U1505 ( .IN1(n1601), .IN2(n1602), .QN(n1604) );
  AO21X1 U1506 ( .IN1(N165), .IN2(n1588), .IN3(n1589), .Q(n1585) );
  XNOR3X1 U1507 ( .IN1(n1605), .IN2(n1606), .IN3(n1607), .Q(n1583) );
  XNOR3X1 U1508 ( .IN1(n1608), .IN2(n1609), .IN3(n1610), .Q(n1607) );
  NAND2X0 U1509 ( .IN1(n1611), .IN2(keyinput100), .QN(n1610) );
  MUX21X1 U1510 ( .IN1(n1612), .IN2(n1613), .S(n1614), .Q(n1611) );
  XOR2X1 U1511 ( .IN1(n1615), .IN2(n1616), .Q(n1614) );
  NOR2X0 U1512 ( .IN1(n1617), .IN2(keyinput41), .QN(n1615) );
  XOR2X1 U1513 ( .IN1(n1618), .IN2(n1619), .Q(n1613) );
  XOR2X1 U1514 ( .IN1(n1620), .IN2(n1619), .Q(n1612) );
  XNOR2X1 U1515 ( .IN1(n1621), .IN2(n1622), .Q(n1619) );
  NAND2X0 U1516 ( .IN1(keyinput91), .IN2(n1618), .QN(n1620) );
  AO221X1 U1517 ( .IN1(n1623), .IN2(N18), .IN3(n1624), .IN4(n1625), .IN5(n1626), .Q(n1618) );
  XOR2X1 U1518 ( .IN1(keyinput53), .IN2(n1627), .Q(n1626) );
  NOR2X0 U1519 ( .IN1(n1628), .IN2(n1629), .QN(n1627) );
  MUX21X1 U1520 ( .IN1(n1630), .IN2(n1625), .S(n1119), .Q(n1629) );
  INVX0 U1521 ( .INP(N44), .ZN(n1625) );
  AND2X1 U1522 ( .IN1(n1630), .IN2(n1628), .Q(n1623) );
  INVX0 U1523 ( .INP(N208), .ZN(n1630) );
  XOR2X1 U1524 ( .IN1(n1631), .IN2(n1632), .Q(n1582) );
  XOR3X1 U1525 ( .IN1(n1633), .IN2(n1634), .IN3(n1635), .Q(n1632) );
  XOR2X1 U1526 ( .IN1(n1636), .IN2(n1637), .Q(n1635) );
  OA21X1 U1527 ( .IN1(n1638), .IN2(n1639), .IN3(n1640), .Q(n1637) );
  XOR2X1 U1528 ( .IN1(n1641), .IN2(keyinput54), .Q(n1640) );
  NAND2X0 U1529 ( .IN1(n1638), .IN2(n1639), .QN(n1641) );
  INVX0 U1530 ( .INP(n1642), .ZN(n1638) );
  NOR2X0 U1531 ( .IN1(keyinput44), .IN2(n1643), .QN(n1636) );
  XNOR3X1 U1532 ( .IN1(n1644), .IN2(n1645), .IN3(n1646), .Q(n1631) );
  MUX21X1 U1533 ( .IN1(n1647), .IN2(n1648), .S(n1122), .Q(n1646) );
  XOR2X1 U1534 ( .IN1(N115), .IN2(n1649), .Q(n1648) );
  XOR2X1 U1535 ( .IN1(N197), .IN2(n1649), .Q(n1647) );
  NOR2X0 U1536 ( .IN1(keyinput40), .IN2(n1650), .QN(n1649) );
  INVX0 U1537 ( .INP(n1651), .ZN(n1650) );
  XNOR2X1 U1538 ( .IN1(n1652), .IN2(n1653), .Q(n1645) );
  MUX41X1 U1539 ( .IN1(n1654), .IN3(n1655), .IN2(n1655), .IN4(n1654), .S0(
        n1656), .S1(n1657), .Q(n1581) );
  AOI21X1 U1540 ( .IN1(N173), .IN2(n1588), .IN3(n1589), .QN(n1657) );
  XOR2X1 U1541 ( .IN1(n1654), .IN2(keyinput74), .Q(n1655) );
  XNOR3X1 U1542 ( .IN1(n1658), .IN2(n1659), .IN3(n1660), .Q(n1654) );
  XNOR3X1 U1543 ( .IN1(n1661), .IN2(n1662), .IN3(n1663), .Q(n1660) );
  XNOR3X1 U1544 ( .IN1(n1664), .IN2(n1665), .IN3(n1666), .Q(n1659) );
  MUX21X1 U1545 ( .IN1(n1667), .IN2(n1668), .S(n1121), .Q(n1666) );
  MUX21X1 U1546 ( .IN1(n1669), .IN2(n1670), .S(N141), .Q(n1668) );
  MUX21X1 U1547 ( .IN1(n1669), .IN2(n1670), .S(N181), .Q(n1667) );
  XNOR2X1 U1548 ( .IN1(n1669), .IN2(keyinput42), .Q(n1670) );
  XNOR2X1 U1549 ( .IN1(n1671), .IN2(n1672), .Q(n1664) );
  XOR2X1 U1550 ( .IN1(keyinput99), .IN2(keyinput59), .Q(n1658) );
  NAND4X0 U1551 ( .IN1(n1673), .IN2(n1674), .IN3(n1675), .IN4(n1676), .QN(
        N10575) );
  XNOR3X1 U1552 ( .IN1(n1677), .IN2(n1678), .IN3(n1679), .Q(n1676) );
  XNOR3X1 U1553 ( .IN1(n1680), .IN2(n1681), .IN3(n1682), .Q(n1679) );
  NAND2X0 U1554 ( .IN1(n1683), .IN2(n1684), .QN(n1682) );
  XNOR2X1 U1555 ( .IN1(n1685), .IN2(keyinput96), .Q(n1684) );
  NAND3X0 U1556 ( .IN1(n1686), .IN2(n1687), .IN3(n1688), .QN(n1685) );
  XNOR2X1 U1557 ( .IN1(n1689), .IN2(keyinput92), .Q(n1688) );
  INVX0 U1558 ( .INP(n1690), .ZN(n1686) );
  MUX21X1 U1559 ( .IN1(n1691), .IN2(n1692), .S(n1690), .Q(n1683) );
  MUX21X1 U1560 ( .IN1(n1693), .IN2(n1694), .S(n1120), .Q(n1690) );
  XNOR2X1 U1561 ( .IN1(N70), .IN2(n1695), .Q(n1694) );
  XOR2X1 U1562 ( .IN1(n1695), .IN2(N310), .Q(n1693) );
  MUX21X1 U1563 ( .IN1(N307), .IN2(n1696), .S(n1119), .Q(n1695) );
  INVX0 U1564 ( .INP(N69), .ZN(n1696) );
  XNOR2X1 U1565 ( .IN1(n1697), .IN2(n1689), .Q(n1692) );
  NAND2X0 U1566 ( .IN1(n1697), .IN2(n1689), .QN(n1691) );
  XNOR2X1 U1567 ( .IN1(n1698), .IN2(n1699), .Q(n1689) );
  INVX0 U1568 ( .INP(n1687), .ZN(n1697) );
  AO21X1 U1569 ( .IN1(n1700), .IN2(n1701), .IN3(n1702), .Q(n1687) );
  XOR2X1 U1570 ( .IN1(keyinput65), .IN2(n1703), .Q(n1702) );
  NOR2X0 U1571 ( .IN1(n1700), .IN2(n1701), .QN(n1703) );
  XOR3X1 U1572 ( .IN1(n1704), .IN2(n1705), .IN3(n1706), .Q(n1675) );
  XNOR3X1 U1573 ( .IN1(n1707), .IN2(n1708), .IN3(n1709), .Q(n1706) );
  MUX21X1 U1574 ( .IN1(n1710), .IN2(n1711), .S(n1122), .Q(n1709) );
  XNOR2X1 U1575 ( .IN1(N114), .IN2(n1712), .Q(n1711) );
  XNOR2X1 U1576 ( .IN1(n1713), .IN2(N248), .Q(n1710) );
  MUX21X1 U1577 ( .IN1(N263), .IN2(n1714), .S(n1121), .Q(n1705) );
  XOR2X1 U1578 ( .IN1(n1715), .IN2(n1716), .Q(n1704) );
  MUX21X1 U1579 ( .IN1(N267), .IN2(n1717), .S(n1120), .Q(n1716) );
  OA21X1 U1580 ( .IN1(n1718), .IN2(n1719), .IN3(n1720), .Q(n1715) );
  XOR2X1 U1581 ( .IN1(n1721), .IN2(keyinput52), .Q(n1720) );
  NAND2X0 U1582 ( .IN1(n1722), .IN2(n1718), .QN(n1721) );
  XOR2X1 U1583 ( .IN1(n1719), .IN2(keyinput38), .Q(n1722) );
  XOR2X1 U1584 ( .IN1(n1723), .IN2(n1724), .Q(n1674) );
  XNOR3X1 U1585 ( .IN1(n1725), .IN2(n1726), .IN3(n1727), .Q(n1724) );
  XNOR3X1 U1586 ( .IN1(keyinput62), .IN2(n1728), .IN3(n1729), .Q(n1723) );
  NAND2X0 U1587 ( .IN1(n1730), .IN2(n1731), .QN(n1729) );
  XOR2X1 U1588 ( .IN1(n1732), .IN2(keyinput86), .Q(n1731) );
  NAND3X0 U1589 ( .IN1(n1733), .IN2(n1734), .IN3(n1735), .QN(n1732) );
  MUX21X1 U1590 ( .IN1(n1736), .IN2(n1737), .S(n1733), .Q(n1730) );
  XOR2X1 U1591 ( .IN1(n1738), .IN2(n1739), .Q(n1733) );
  NAND2X0 U1592 ( .IN1(keyinput43), .IN2(n1740), .QN(n1738) );
  OR2X1 U1593 ( .IN1(n1735), .IN2(n1734), .Q(n1737) );
  XNOR2X1 U1594 ( .IN1(n1734), .IN2(n1735), .Q(n1736) );
  XOR3X1 U1595 ( .IN1(keyinput60), .IN2(n1741), .IN3(n1742), .Q(n1735) );
  MUX21X1 U1596 ( .IN1(n1743), .IN2(N82), .S(n1119), .Q(n1741) );
  INVX0 U1597 ( .INP(N274), .ZN(n1743) );
  XOR2X1 U1598 ( .IN1(n1744), .IN2(n1745), .Q(n1734) );
  XNOR3X1 U1599 ( .IN1(n1746), .IN2(n1747), .IN3(n1748), .Q(n1673) );
  XOR2X1 U1600 ( .IN1(n1749), .IN2(n1750), .Q(n1748) );
  NOR2X0 U1601 ( .IN1(keyinput107), .IN2(n1751), .QN(n1750) );
  XOR3X1 U1602 ( .IN1(n1752), .IN2(n1753), .IN3(n1754), .Q(n1751) );
  OA21X1 U1603 ( .IN1(n1755), .IN2(n1756), .IN3(n1757), .Q(n1752) );
  XOR2X1 U1604 ( .IN1(n1758), .IN2(keyinput66), .Q(n1757) );
  NAND2X0 U1605 ( .IN1(n1755), .IN2(n1756), .QN(n1758) );
  NAND2X0 U1606 ( .IN1(keyinput80), .IN2(n1759), .QN(n1749) );
  XNOR3X1 U1607 ( .IN1(n1760), .IN2(n1761), .IN3(n1762), .Q(n1759) );
  MUX21X1 U1608 ( .IN1(n1763), .IN2(n1764), .S(n1122), .Q(n1762) );
  XNOR2X1 U1609 ( .IN1(n1765), .IN2(N58), .Q(n1764) );
  XOR2X1 U1610 ( .IN1(N337), .IN2(n1765), .Q(n1763) );
  NAND4X0 U1611 ( .IN1(n1766), .IN2(n1767), .IN3(n1768), .IN4(n1769), .QN(
        N10574) );
  XOR3X1 U1612 ( .IN1(n1770), .IN2(n1771), .IN3(n1772), .Q(n1769) );
  XOR3X1 U1613 ( .IN1(n1773), .IN2(n1546), .IN3(n1774), .Q(n1772) );
  AOI21X1 U1614 ( .IN1(n1775), .IN2(keyinput77), .IN3(n1776), .QN(n1774) );
  INVX0 U1615 ( .INP(n1777), .ZN(n1776) );
  MUX21X1 U1616 ( .IN1(n1778), .IN2(n1779), .S(n1780), .Q(n1777) );
  XNOR2X1 U1617 ( .IN1(n1781), .IN2(n1782), .Q(n1780) );
  NAND2X0 U1618 ( .IN1(keyinput29), .IN2(n1544), .QN(n1781) );
  OA22X1 U1619 ( .IN1(keyinput77), .IN2(n1775), .IN3(n1783), .IN4(n1784), .Q(
        n1779) );
  NOR2X0 U1620 ( .IN1(keyinput77), .IN2(n1785), .QN(n1778) );
  XNOR2X1 U1621 ( .IN1(n1786), .IN2(n1784), .Q(n1785) );
  NAND2X0 U1622 ( .IN1(keyinput76), .IN2(n1783), .QN(n1786) );
  NAND2X0 U1623 ( .IN1(n1783), .IN2(n1784), .QN(n1775) );
  XNOR2X1 U1624 ( .IN1(n1787), .IN2(n1788), .Q(n1784) );
  MUX21X1 U1625 ( .IN1(n1789), .IN2(n1790), .S(n1121), .Q(n1783) );
  XNOR2X1 U1626 ( .IN1(n1384), .IN2(N141), .Q(n1790) );
  XNOR2X1 U1627 ( .IN1(n1384), .IN2(N161), .Q(n1789) );
  XNOR2X1 U1628 ( .IN1(n1791), .IN2(n1548), .Q(n1771) );
  XOR2X1 U1629 ( .IN1(keyinput97), .IN2(keyinput61), .Q(n1770) );
  XOR2X1 U1630 ( .IN1(n1792), .IN2(n1793), .Q(n1768) );
  XNOR3X1 U1631 ( .IN1(n1503), .IN2(n1794), .IN3(n1795), .Q(n1793) );
  XNOR2X1 U1632 ( .IN1(n1796), .IN2(n1797), .Q(n1795) );
  XOR3X1 U1633 ( .IN1(n1798), .IN2(n1799), .IN3(n1800), .Q(n1792) );
  AO21X1 U1634 ( .IN1(N211), .IN2(n1801), .IN3(n1802), .Q(n1800) );
  AO21X1 U1635 ( .IN1(N212), .IN2(n1801), .IN3(n1802), .Q(n1799) );
  NAND2X0 U1636 ( .IN1(n1803), .IN2(n1801), .QN(n1798) );
  XNOR3X1 U1637 ( .IN1(n1804), .IN2(n1805), .IN3(n1806), .Q(n1767) );
  XOR2X1 U1638 ( .IN1(n1807), .IN2(n1808), .Q(n1806) );
  XNOR3X1 U1639 ( .IN1(keyinput71), .IN2(n1809), .IN3(n1810), .Q(n1808) );
  XNOR2X1 U1640 ( .IN1(n1811), .IN2(n1812), .Q(n1810) );
  XNOR3X1 U1641 ( .IN1(n1533), .IN2(n1813), .IN3(n1814), .Q(n1807) );
  MUX21X1 U1642 ( .IN1(n1815), .IN2(n1816), .S(n1120), .Q(n1814) );
  XNOR2X1 U1643 ( .IN1(N44), .IN2(n1817), .Q(n1816) );
  XNOR2X1 U1644 ( .IN1(N239), .IN2(n1817), .Q(n1815) );
  XNOR2X1 U1645 ( .IN1(n1818), .IN2(n1819), .Q(n1813) );
  XNOR3X1 U1646 ( .IN1(n1820), .IN2(n1821), .IN3(n1822), .Q(n1766) );
  XOR3X1 U1647 ( .IN1(n1515), .IN2(n1823), .IN3(n1824), .Q(n1822) );
  MUX21X1 U1648 ( .IN1(n1825), .IN2(n1826), .S(n1119), .Q(n1824) );
  XOR2X1 U1649 ( .IN1(N115), .IN2(n1827), .Q(n1826) );
  XOR2X1 U1650 ( .IN1(N227), .IN2(n1827), .Q(n1825) );
  XNOR2X1 U1651 ( .IN1(n1828), .IN2(n1829), .Q(n1823) );
  XNOR3X1 U1652 ( .IN1(n1537), .IN2(n1830), .IN3(n1831), .Q(n1820) );
  XNOR2X1 U1653 ( .IN1(n1832), .IN2(n1833), .Q(n1831) );
  XNOR3X1 U1654 ( .IN1(keyinput111), .IN2(n1430), .IN3(n1834), .Q(N10353) );
  MUX21X1 U1655 ( .IN1(n1835), .IN2(n1836), .S(n1430), .Q(N10352) );
  XNOR2X1 U1656 ( .IN1(n1179), .IN2(n1523), .Q(n1836) );
  AO21X1 U1657 ( .IN1(n1837), .IN2(n1523), .IN3(n1838), .Q(n1835) );
  XOR2X1 U1658 ( .IN1(keyinput94), .IN2(n1839), .Q(n1838) );
  NOR2X0 U1659 ( .IN1(n1523), .IN2(n1837), .QN(n1839) );
  INVX0 U1660 ( .INP(n1183), .ZN(n1523) );
  MUX21X1 U1661 ( .IN1(n1840), .IN2(n1841), .S(n1430), .Q(N10351) );
  XNOR2X1 U1662 ( .IN1(n1842), .IN2(n1174), .Q(n1841) );
  AOI21X1 U1663 ( .IN1(n1161), .IN2(n1843), .IN3(n1844), .QN(n1840) );
  MUX21X1 U1664 ( .IN1(n1845), .IN2(n1846), .S(n1430), .Q(N10350) );
  XNOR2X1 U1665 ( .IN1(n1184), .IN2(n1847), .Q(n1846) );
  OA21X1 U1666 ( .IN1(n1842), .IN2(n1161), .IN3(n1848), .Q(n1847) );
  INVX0 U1667 ( .INP(n1522), .ZN(n1848) );
  NOR2X0 U1668 ( .IN1(n1849), .IN2(n1175), .QN(n1842) );
  INVX0 U1669 ( .INP(n1843), .ZN(n1849) );
  NOR2X0 U1670 ( .IN1(n1850), .IN2(n1851), .QN(n1845) );
  NOR3X0 U1671 ( .IN1(n1844), .IN2(n1184), .IN3(n1522), .QN(n1851) );
  XOR2X1 U1672 ( .IN1(n1159), .IN2(n1852), .Q(N10112) );
  XNOR2X1 U1673 ( .IN1(n1158), .IN2(n1853), .Q(N10111) );
  XNOR2X1 U1674 ( .IN1(n1854), .IN2(n1855), .Q(N10110) );
  NOR2X0 U1675 ( .IN1(n1856), .IN2(n1857), .QN(n1855) );
  XNOR2X1 U1676 ( .IN1(n1141), .IN2(n1858), .Q(N10109) );
  OA21X1 U1677 ( .IN1(n1859), .IN2(n1860), .IN3(n1528), .Q(n1858) );
  INVX0 U1678 ( .INP(n1861), .ZN(n1528) );
  INVX0 U1679 ( .INP(n1854), .ZN(n1860) );
  OA21X1 U1680 ( .IN1(n1853), .IN2(n1529), .IN3(n1530), .Q(n1859) );
  INVX0 U1681 ( .INP(n1862), .ZN(n1530) );
  OA21X1 U1682 ( .IN1(n1159), .IN2(n1852), .IN3(n1863), .Q(n1853) );
  OA21X1 U1683 ( .IN1(n1128), .IN2(n1131), .IN3(n1138), .Q(n1852) );
  NAND3X0 U1684 ( .IN1(n1864), .IN2(n1865), .IN3(n1574), .QN(N10102) );
  OA21X1 U1685 ( .IN1(n1866), .IN2(n1867), .IN3(n1868), .Q(n1574) );
  XNOR2X1 U1686 ( .IN1(n1869), .IN2(keyinput8), .Q(n1868) );
  NAND2X0 U1687 ( .IN1(N38), .IN2(n1867), .QN(n1869) );
  OR2X1 U1688 ( .IN1(n1578), .IN2(n1580), .Q(n1865) );
  NAND4X0 U1689 ( .IN1(n1870), .IN2(n1871), .IN3(n1872), .IN4(n1873), .QN(
        n1578) );
  NOR3X0 U1690 ( .IN1(n1874), .IN2(n1875), .IN3(n1876), .QN(n1873) );
  XNOR2X1 U1691 ( .IN1(n1600), .IN2(n1712), .Q(n1874) );
  INVX0 U1692 ( .INP(n1713), .ZN(n1712) );
  NAND2X0 U1693 ( .IN1(n1877), .IN2(n1878), .QN(n1871) );
  AO221X1 U1694 ( .IN1(n1879), .IN2(n1880), .IN3(n1728), .IN4(n1656), .IN5(
        n1881), .Q(n1878) );
  XNOR2X1 U1695 ( .IN1(n1882), .IN2(n1883), .Q(n1881) );
  OA21X1 U1696 ( .IN1(n1661), .IN2(n1884), .IN3(n1885), .Q(n1880) );
  OAI221X1 U1697 ( .IN1(n1886), .IN2(n1887), .IN3(n1888), .IN4(n1662), .IN5(
        n1889), .QN(n1885) );
  AND2X1 U1698 ( .IN1(n1662), .IN2(n1888), .Q(n1887) );
  AO21X1 U1699 ( .IN1(n1739), .IN2(n1663), .IN3(n1890), .Q(n1888) );
  OA221X1 U1700 ( .IN1(n1891), .IN2(n1671), .IN3(n1892), .IN4(n1740), .IN5(
        n1893), .Q(n1890) );
  AND2X1 U1701 ( .IN1(n1671), .IN2(n1891), .Q(n1892) );
  AOI22X1 U1702 ( .IN1(n1665), .IN2(n1894), .IN3(n1745), .IN4(n1895), .QN(
        n1891) );
  OR2X1 U1703 ( .IN1(n1894), .IN2(n1665), .Q(n1895) );
  INVX0 U1704 ( .INP(n1896), .ZN(n1745) );
  AO22X1 U1705 ( .IN1(n1897), .IN2(n1898), .IN3(n1744), .IN4(n1899), .Q(n1894)
         );
  OR2X1 U1706 ( .IN1(n1897), .IN2(n1898), .Q(n1899) );
  INVX0 U1707 ( .INP(n1900), .ZN(n1744) );
  INVX0 U1708 ( .INP(n1672), .ZN(n1898) );
  XNOR2X1 U1709 ( .IN1(n1901), .IN2(keyinput25), .Q(n1897) );
  NAND2X0 U1710 ( .IN1(n1742), .IN2(n1902), .QN(n1901) );
  INVX0 U1711 ( .INP(n1903), .ZN(n1665) );
  OA21X1 U1712 ( .IN1(n1728), .IN2(n1656), .IN3(n1904), .Q(n1879) );
  NAND4X0 U1713 ( .IN1(n1905), .IN2(n1889), .IN3(n1906), .IN4(n1907), .QN(
        n1904) );
  OA221X1 U1714 ( .IN1(n1672), .IN2(n1900), .IN3(n1903), .IN4(n1896), .IN5(
        n1908), .Q(n1907) );
  OA21X1 U1715 ( .IN1(n1662), .IN2(n1886), .IN3(n1893), .Q(n1908) );
  MUX21X1 U1716 ( .IN1(n1909), .IN2(n1910), .S(keyinput56), .Q(n1893) );
  NOR2X0 U1717 ( .IN1(n1663), .IN2(n1739), .QN(n1910) );
  OR2X1 U1718 ( .IN1(n1739), .IN2(n1663), .Q(n1909) );
  OA21X1 U1719 ( .IN1(N177), .IN2(n1589), .IN3(n1588), .Q(n1663) );
  MUX21X1 U1720 ( .IN1(n1911), .IN2(N64), .S(n1122), .Q(n1739) );
  INVX0 U1721 ( .INP(N289), .ZN(n1911) );
  INVX0 U1722 ( .INP(n1726), .ZN(n1886) );
  MUX21X1 U1723 ( .IN1(N293), .IN2(n1912), .S(n1121), .Q(n1726) );
  INVX0 U1724 ( .INP(N63), .ZN(n1912) );
  AO21X1 U1725 ( .IN1(N176), .IN2(n1588), .IN3(n1589), .Q(n1662) );
  MUX21X1 U1726 ( .IN1(n1541), .IN2(N84), .S(n1120), .Q(n1896) );
  MUX21X1 U1727 ( .IN1(N179), .IN2(N144), .S(n1119), .Q(n1903) );
  MUX21X1 U1728 ( .IN1(n1913), .IN2(N83), .S(n1122), .Q(n1900) );
  MUX21X1 U1729 ( .IN1(N180), .IN2(N138), .S(n1121), .Q(n1672) );
  OA22X1 U1730 ( .IN1(n1914), .IN2(n1915), .IN3(n1671), .IN4(n1740), .Q(n1906)
         );
  AO21X1 U1731 ( .IN1(N85), .IN2(n1121), .IN3(n1916), .Q(n1740) );
  XOR2X1 U1732 ( .IN1(keyinput15), .IN2(n1917), .Q(n1916) );
  NOR2X0 U1733 ( .IN1(N286), .IN2(n1122), .QN(n1917) );
  MUX21X1 U1734 ( .IN1(N178), .IN2(N135), .S(n1120), .Q(n1671) );
  XOR2X1 U1735 ( .IN1(n1918), .IN2(keyinput48), .Q(n1915) );
  NAND2X0 U1736 ( .IN1(n1742), .IN2(n1669), .QN(n1918) );
  NOR2X0 U1737 ( .IN1(n1669), .IN2(n1742), .QN(n1914) );
  MUX21X1 U1738 ( .IN1(n1919), .IN2(N65), .S(n1119), .Q(n1742) );
  INVX0 U1739 ( .INP(n1902), .ZN(n1669) );
  MUX21X1 U1740 ( .IN1(N171), .IN2(N147), .S(n1122), .Q(n1902) );
  NAND2X0 U1741 ( .IN1(n1884), .IN2(n1661), .QN(n1889) );
  OAI21X1 U1742 ( .IN1(N175), .IN2(n1589), .IN3(n1588), .QN(n1661) );
  INVX0 U1743 ( .INP(n1725), .ZN(n1884) );
  MUX21X1 U1744 ( .IN1(n1920), .IN2(N86), .S(n1121), .Q(n1725) );
  AO221X1 U1745 ( .IN1(n1921), .IN2(n1554), .IN3(n1922), .IN4(n1923), .IN5(
        n1557), .Q(n1905) );
  AO22X1 U1746 ( .IN1(n1634), .IN2(n1753), .IN3(n1924), .IN4(n1925), .Q(n1557)
         );
  AO22X1 U1747 ( .IN1(n1754), .IN2(n1926), .IN3(n1927), .IN4(n1928), .Q(n1925)
         );
  NAND2X0 U1748 ( .IN1(n1929), .IN2(n1930), .QN(n1928) );
  NAND3X0 U1749 ( .IN1(n1756), .IN2(n1642), .IN3(n1931), .QN(n1929) );
  INVX0 U1750 ( .INP(n1932), .ZN(n1756) );
  AND3X1 U1751 ( .IN1(n1563), .IN2(n1565), .IN3(n1933), .Q(n1923) );
  OAI21X1 U1752 ( .IN1(n1570), .IN2(n1569), .IN3(n1934), .QN(n1933) );
  XNOR2X1 U1753 ( .IN1(keyinput101), .IN2(n1935), .Q(n1934) );
  OA21X1 U1754 ( .IN1(n1568), .IN2(n1570), .IN3(n1566), .Q(n1935) );
  XOR2X1 U1755 ( .IN1(keyinput85), .IN2(n1936), .Q(n1566) );
  OA21X1 U1756 ( .IN1(n1937), .IN2(n1938), .IN3(n1939), .Q(n1936) );
  OA22X1 U1757 ( .IN1(n1940), .IN2(n1941), .IN3(n1942), .IN4(n1677), .Q(n1937)
         );
  INVX0 U1758 ( .INP(n1943), .ZN(n1941) );
  OA21X1 U1759 ( .IN1(n1605), .IN2(n1681), .IN3(n1944), .Q(n1940) );
  NAND3X0 U1760 ( .IN1(n1945), .IN2(n1608), .IN3(n1678), .QN(n1944) );
  INVX0 U1761 ( .INP(n1946), .ZN(n1605) );
  AOI221X1 U1762 ( .IN1(n1947), .IN2(n1622), .IN3(n1948), .IN4(n1949), .IN5(
        n1950), .QN(n1568) );
  XNOR2X1 U1763 ( .IN1(n1951), .IN2(keyinput79), .Q(n1950) );
  NAND3X0 U1764 ( .IN1(n1624), .IN2(n1952), .IN3(n1953), .QN(n1951) );
  AO22X1 U1765 ( .IN1(n1698), .IN2(n1621), .IN3(n1954), .IN4(n1955), .Q(n1949)
         );
  AO22X1 U1766 ( .IN1(n1956), .IN2(n1616), .IN3(n1957), .IN4(n1958), .Q(n1955)
         );
  NOR2X0 U1767 ( .IN1(n1617), .IN2(n1959), .QN(n1957) );
  INVX0 U1768 ( .INP(n1700), .ZN(n1956) );
  INVX0 U1769 ( .INP(n1960), .ZN(n1698) );
  INVX0 U1770 ( .INP(n1699), .ZN(n1947) );
  NAND3X0 U1771 ( .IN1(n1953), .IN2(n1961), .IN3(N89), .QN(n1569) );
  XOR2X1 U1772 ( .IN1(n1624), .IN2(n1952), .Q(n1961) );
  XNOR2X1 U1773 ( .IN1(n1962), .IN2(keyinput20), .Q(n1952) );
  OR2X1 U1774 ( .IN1(N70), .IN2(N18), .Q(n1962) );
  AND2X1 U1775 ( .IN1(n1628), .IN2(n1122), .Q(n1624) );
  MUX21X1 U1776 ( .IN1(N198), .IN2(N41), .S(n1120), .Q(n1628) );
  AND4X1 U1777 ( .IN1(n1963), .IN2(n1958), .IN3(n1954), .IN4(n1948), .Q(n1953)
         );
  XNOR2X1 U1778 ( .IN1(n1699), .IN2(n1622), .Q(n1948) );
  MUX21X1 U1779 ( .IN1(N204), .IN2(N103), .S(n1119), .Q(n1622) );
  MUX21X1 U1780 ( .IN1(N322), .IN2(n1964), .S(n1122), .Q(n1699) );
  INVX0 U1781 ( .INP(N73), .ZN(n1964) );
  XNOR2X1 U1782 ( .IN1(n1960), .IN2(n1621), .Q(n1954) );
  MUX21X1 U1783 ( .IN1(N205), .IN2(N23), .S(n1121), .Q(n1621) );
  MUX21X1 U1784 ( .IN1(N319), .IN2(n1965), .S(n1120), .Q(n1960) );
  INVX0 U1785 ( .INP(N75), .ZN(n1965) );
  XNOR2X1 U1786 ( .IN1(n1700), .IN2(n1616), .Q(n1958) );
  MUX21X1 U1787 ( .IN1(N206), .IN2(N26), .S(n1119), .Q(n1616) );
  MUX21X1 U1788 ( .IN1(n1966), .IN2(n1967), .S(n1122), .Q(n1700) );
  INVX0 U1789 ( .INP(N76), .ZN(n1967) );
  XNOR2X1 U1790 ( .IN1(n1701), .IN2(n1617), .Q(n1963) );
  AOI21X1 U1791 ( .IN1(N29), .IN2(n1120), .IN3(n1968), .QN(n1617) );
  XNOR2X1 U1792 ( .IN1(n1969), .IN2(keyinput16), .Q(n1968) );
  NAND2X0 U1793 ( .IN1(N207), .IN2(N18), .QN(n1969) );
  INVX0 U1794 ( .INP(n1959), .ZN(n1701) );
  MUX21X1 U1795 ( .IN1(N313), .IN2(n1970), .S(n1121), .Q(n1959) );
  INVX0 U1796 ( .INP(N74), .ZN(n1970) );
  NAND4X0 U1797 ( .IN1(n1971), .IN2(n1972), .IN3(n1943), .IN4(n1945), .QN(
        n1570) );
  AO21X1 U1798 ( .IN1(n1681), .IN2(n1946), .IN3(n1973), .Q(n1945) );
  XOR2X1 U1799 ( .IN1(keyinput64), .IN2(n1974), .Q(n1973) );
  NOR2X0 U1800 ( .IN1(n1946), .IN2(n1681), .QN(n1974) );
  MUX21X1 U1801 ( .IN1(N202), .IN2(N127), .S(n1120), .Q(n1946) );
  MUX21X1 U1802 ( .IN1(n1975), .IN2(n1976), .S(N18), .Q(n1681) );
  INVX0 U1803 ( .INP(N54), .ZN(n1975) );
  XOR2X1 U1804 ( .IN1(n1677), .IN2(n1942), .Q(n1943) );
  INVX0 U1805 ( .INP(n1606), .ZN(n1942) );
  MUX21X1 U1806 ( .IN1(N201), .IN2(N124), .S(n1119), .Q(n1606) );
  MUX21X1 U1807 ( .IN1(N331), .IN2(n1977), .S(n1122), .Q(n1677) );
  INVX0 U1808 ( .INP(N55), .ZN(n1977) );
  INVX0 U1809 ( .INP(n1938), .ZN(n1972) );
  MUX21X1 U1810 ( .IN1(n1978), .IN2(n1979), .S(keyinput72), .Q(n1938) );
  OA21X1 U1811 ( .IN1(n1680), .IN2(n1609), .IN3(n1939), .Q(n1979) );
  NAND2X0 U1812 ( .IN1(n1680), .IN2(n1609), .QN(n1939) );
  XNOR2X1 U1813 ( .IN1(n1680), .IN2(n1609), .Q(n1978) );
  XNOR2X1 U1814 ( .IN1(n1980), .IN2(keyinput23), .Q(n1609) );
  MUX21X1 U1815 ( .IN1(N200), .IN2(N100), .S(n1121), .Q(n1980) );
  MUX21X1 U1816 ( .IN1(n1981), .IN2(N56), .S(n1120), .Q(n1680) );
  XOR2X1 U1817 ( .IN1(n1678), .IN2(n1608), .Q(n1971) );
  AO21X1 U1818 ( .IN1(N130), .IN2(n1119), .IN3(n1982), .Q(n1608) );
  XOR2X1 U1819 ( .IN1(n1983), .IN2(keyinput21), .Q(n1982) );
  NAND2X0 U1820 ( .IN1(N203), .IN2(N18), .QN(n1983) );
  MUX21X1 U1821 ( .IN1(n1984), .IN2(N53), .S(n1119), .Q(n1678) );
  OA22X1 U1822 ( .IN1(n1760), .IN2(n1985), .IN3(n1651), .IN4(n1765), .Q(n1563)
         );
  AND2X1 U1823 ( .IN1(n1562), .IN2(n1554), .Q(n1922) );
  AND4X1 U1824 ( .IN1(n1924), .IN2(n1931), .IN3(n1986), .IN4(n1927), .Q(n1554)
         );
  XNOR2X1 U1825 ( .IN1(n1643), .IN2(n1754), .Q(n1927) );
  MUX21X1 U1826 ( .IN1(n1987), .IN2(N61), .S(n1122), .Q(n1754) );
  INVX0 U1827 ( .INP(n1926), .ZN(n1643) );
  MUX21X1 U1828 ( .IN1(N190), .IN2(N50), .S(n1121), .Q(n1926) );
  XNOR2X1 U1829 ( .IN1(n1642), .IN2(n1932), .Q(n1986) );
  MUX21X1 U1830 ( .IN1(N355), .IN2(n1988), .S(n1120), .Q(n1932) );
  INVX0 U1831 ( .INP(N79), .ZN(n1988) );
  MUX21X1 U1832 ( .IN1(N192), .IN2(N35), .S(n1119), .Q(n1642) );
  AOI22X1 U1833 ( .IN1(n1989), .IN2(keyinput57), .IN3(n1755), .IN4(n1990), 
        .QN(n1931) );
  NAND2X0 U1834 ( .IN1(keyinput57), .IN2(n1639), .QN(n1990) );
  INVX0 U1835 ( .INP(n1991), .ZN(n1755) );
  INVX0 U1836 ( .INP(n1930), .ZN(n1989) );
  NAND2X0 U1837 ( .IN1(n1991), .IN2(n1639), .QN(n1930) );
  MUX21X1 U1838 ( .IN1(N32), .IN2(N191), .S(N18), .Q(n1639) );
  MUX21X1 U1839 ( .IN1(n1992), .IN2(N60), .S(n1122), .Q(n1991) );
  XOR2X1 U1840 ( .IN1(n1753), .IN2(n1634), .Q(n1924) );
  MUX21X1 U1841 ( .IN1(N189), .IN2(N66), .S(n1121), .Q(n1634) );
  AO21X1 U1842 ( .IN1(N18), .IN2(n1516), .IN3(n1993), .Q(n1753) );
  XOR2X1 U1843 ( .IN1(n1994), .IN2(keyinput17), .Q(n1993) );
  NAND2X0 U1844 ( .IN1(N62), .IN2(n1121), .QN(n1994) );
  INVX0 U1845 ( .INP(n1560), .ZN(n1921) );
  AO22X1 U1846 ( .IN1(n1995), .IN2(n1996), .IN3(n1653), .IN4(n1997), .Q(n1560)
         );
  OR2X1 U1847 ( .IN1(n1996), .IN2(n1995), .Q(n1997) );
  INVX0 U1848 ( .INP(n1985), .ZN(n1653) );
  MUX21X1 U1849 ( .IN1(N193), .IN2(N47), .S(n1120), .Q(n1985) );
  NAND2X0 U1850 ( .IN1(n1565), .IN2(n1998), .QN(n1996) );
  AO221X1 U1851 ( .IN1(n1562), .IN2(n1999), .IN3(n1761), .IN4(n1633), .IN5(
        n2000), .Q(n1998) );
  XOR2X1 U1852 ( .IN1(n2001), .IN2(keyinput36), .Q(n2000) );
  NAND2X0 U1853 ( .IN1(n1652), .IN2(n1747), .QN(n2001) );
  AO22X1 U1854 ( .IN1(n1765), .IN2(n1651), .IN3(n1746), .IN4(n1644), .Q(n1999)
         );
  MUX21X1 U1855 ( .IN1(N187), .IN2(N118), .S(n1119), .Q(n1651) );
  MUX21X1 U1856 ( .IN1(n2002), .IN2(N77), .S(n1122), .Q(n1765) );
  OA21X1 U1857 ( .IN1(n1746), .IN2(n1644), .IN3(n2003), .Q(n1562) );
  XOR2X1 U1858 ( .IN1(n1652), .IN2(n1747), .Q(n2003) );
  MUX21X1 U1859 ( .IN1(N59), .IN2(n2004), .S(N18), .Q(n1747) );
  MUX21X1 U1860 ( .IN1(N195), .IN2(N94), .S(n1121), .Q(n1652) );
  MUX21X1 U1861 ( .IN1(N196), .IN2(N97), .S(n1120), .Q(n1644) );
  MUX21X1 U1862 ( .IN1(n2005), .IN2(N78), .S(n1119), .Q(n1746) );
  OR2X1 U1863 ( .IN1(n1761), .IN2(n1633), .Q(n1565) );
  MUX21X1 U1864 ( .IN1(N194), .IN2(N121), .S(n1122), .Q(n1633) );
  MUX21X1 U1865 ( .IN1(N81), .IN2(n2006), .S(N18), .Q(n1761) );
  INVX0 U1866 ( .INP(n1760), .ZN(n1995) );
  AO21X1 U1867 ( .IN1(N80), .IN2(n1120), .IN3(n2007), .Q(n1760) );
  XOR2X1 U1868 ( .IN1(n2008), .IN2(keyinput22), .Q(n2007) );
  OR2X1 U1869 ( .IN1(n1121), .IN2(N352), .Q(n2008) );
  AO21X1 U1870 ( .IN1(n2009), .IN2(N18), .IN3(n1600), .Q(n1656) );
  XNOR2X1 U1871 ( .IN1(keyinput9), .IN2(N174), .Q(n2009) );
  MUX21X1 U1872 ( .IN1(N299), .IN2(n2010), .S(n1121), .Q(n1728) );
  INVX0 U1873 ( .INP(N109), .ZN(n2010) );
  XOR2X1 U1874 ( .IN1(n2011), .IN2(keyinput24), .Q(n1877) );
  NAND2X0 U1875 ( .IN1(n1883), .IN2(n1882), .QN(n2011) );
  AO21X1 U1876 ( .IN1(N173), .IN2(n1588), .IN3(n1589), .Q(n1882) );
  INVX0 U1877 ( .INP(n1727), .ZN(n1883) );
  MUX21X1 U1878 ( .IN1(N303), .IN2(n2012), .S(n1120), .Q(n1727) );
  INVX0 U1879 ( .INP(N110), .ZN(n2012) );
  XOR2X1 U1880 ( .IN1(keyinput84), .IN2(n2013), .Q(n1864) );
  NOR2X0 U1881 ( .IN1(n1579), .IN2(n1580), .QN(n2013) );
  NAND2X0 U1882 ( .IN1(n2014), .IN2(n1866), .QN(n1580) );
  NAND2X0 U1883 ( .IN1(N38), .IN2(n2015), .QN(n1866) );
  MUX21X1 U1884 ( .IN1(n2016), .IN2(n2017), .S(n2018), .Q(n2014) );
  AND2X1 U1885 ( .IN1(n1867), .IN2(n2015), .Q(n2017) );
  XNOR2X1 U1886 ( .IN1(n2019), .IN2(keyinput7), .Q(n2015) );
  NAND2X0 U1887 ( .IN1(N382), .IN2(n1714), .QN(n2019) );
  INVX0 U1888 ( .INP(N245), .ZN(n1714) );
  INVX0 U1889 ( .INP(n1867), .ZN(n2016) );
  NAND2X0 U1890 ( .IN1(N382), .IN2(n1717), .QN(n1867) );
  INVX0 U1891 ( .INP(N271), .ZN(n1717) );
  OA22X1 U1892 ( .IN1(n1602), .IN2(n2020), .IN3(n2021), .IN4(n1875), .Q(n1579)
         );
  XNOR2X1 U1893 ( .IN1(n1718), .IN2(n2022), .Q(n1875) );
  OA21X1 U1894 ( .IN1(n2023), .IN2(n1876), .IN3(n2024), .Q(n2021) );
  XOR2X1 U1895 ( .IN1(keyinput26), .IN2(n2025), .Q(n2024) );
  NOR2X0 U1896 ( .IN1(n2026), .IN2(n1719), .QN(n2025) );
  XNOR2X1 U1897 ( .IN1(n2026), .IN2(n1719), .Q(n1876) );
  MUX21X1 U1898 ( .IN1(N257), .IN2(n2027), .S(n1119), .Q(n1719) );
  INVX0 U1899 ( .INP(N112), .ZN(n2027) );
  INVX0 U1900 ( .INP(n1601), .ZN(n2026) );
  AO21X1 U1901 ( .IN1(N167), .IN2(n1588), .IN3(n1589), .Q(n1601) );
  AOI22X1 U1902 ( .IN1(n2028), .IN2(n1870), .IN3(n1599), .IN4(n2029), .QN(
        n2023) );
  AO21X1 U1903 ( .IN1(n1708), .IN2(n1599), .IN3(n2030), .Q(n1870) );
  XOR2X1 U1904 ( .IN1(keyinput49), .IN2(n2031), .Q(n2030) );
  NOR2X0 U1905 ( .IN1(n1599), .IN2(n1708), .QN(n2031) );
  AO21X1 U1906 ( .IN1(N168), .IN2(n1588), .IN3(n1589), .Q(n1599) );
  INVX0 U1907 ( .INP(n2029), .ZN(n1708) );
  MUX21X1 U1908 ( .IN1(n2032), .IN2(N87), .S(n1122), .Q(n2029) );
  OAI21X1 U1909 ( .IN1(n1598), .IN2(n1707), .IN3(n2033), .QN(n2028) );
  NAND3X0 U1910 ( .IN1(n1872), .IN2(n1588), .IN3(n1713), .QN(n2033) );
  XNOR2X1 U1911 ( .IN1(n2034), .IN2(keyinput18), .Q(n1713) );
  MUX21X1 U1912 ( .IN1(n1302), .IN2(N113), .S(n1121), .Q(n2034) );
  AO21X1 U1913 ( .IN1(n1598), .IN2(n2035), .IN3(n2036), .Q(n1872) );
  XOR2X1 U1914 ( .IN1(n2037), .IN2(keyinput50), .Q(n2036) );
  NAND2X0 U1915 ( .IN1(n1707), .IN2(n2038), .QN(n2037) );
  INVX0 U1916 ( .INP(n1707), .ZN(n2035) );
  MUX21X1 U1917 ( .IN1(N254), .IN2(n2039), .S(n1120), .Q(n1707) );
  INVX0 U1918 ( .INP(N111), .ZN(n2039) );
  INVX0 U1919 ( .INP(n2038), .ZN(n1598) );
  AO21X1 U1920 ( .IN1(N169), .IN2(n1588), .IN3(n1589), .Q(n2038) );
  INVX0 U1921 ( .INP(n1718), .ZN(n2020) );
  MUX21X1 U1922 ( .IN1(n2040), .IN2(N88), .S(n1119), .Q(n1718) );
  INVX0 U1923 ( .INP(n2022), .ZN(n1602) );
  OA21X1 U1924 ( .IN1(N166), .IN2(n1589), .IN3(n1588), .Q(n2022) );
  NOR2X0 U1925 ( .IN1(n1600), .IN2(N18), .QN(n1589) );
  INVX0 U1926 ( .INP(n1588), .ZN(n1600) );
  AO21X1 U1927 ( .IN1(n1320), .IN2(n1431), .IN3(n1497), .Q(N10759) );
  AO21X1 U1928 ( .IN1(N38), .IN2(n2041), .IN3(n1433), .Q(n1497) );
  INVX0 U1929 ( .INP(n1317), .ZN(n1433) );
  AO21X1 U1930 ( .IN1(n2042), .IN2(n1471), .IN3(n1499), .Q(n1431) );
  NOR2X0 U1931 ( .IN1(N260), .IN2(n2043), .QN(n1499) );
  NAND2X0 U1932 ( .IN1(n1553), .IN2(n1552), .QN(n1471) );
  NAND2X0 U1933 ( .IN1(n2043), .IN2(n2040), .QN(n1552) );
  INVX0 U1934 ( .INP(N260), .ZN(n2040) );
  INVX0 U1935 ( .INP(n1796), .ZN(n2043) );
  NAND2X0 U1936 ( .IN1(N260), .IN2(n1796), .QN(n1553) );
  AO21X1 U1937 ( .IN1(N213), .IN2(n1801), .IN3(n1802), .Q(n1796) );
  NAND2X0 U1938 ( .IN1(n1311), .IN2(n2044), .QN(n2042) );
  NAND3X0 U1939 ( .IN1(n1469), .IN2(n1468), .IN3(n1295), .QN(n2044) );
  INVX0 U1940 ( .INP(n1306), .ZN(n1295) );
  NAND2X0 U1941 ( .IN1(n1294), .IN2(n2045), .QN(n1468) );
  NAND3X0 U1942 ( .IN1(n1467), .IN2(n1466), .IN3(n1290), .QN(n2045) );
  INVX0 U1943 ( .INP(n1296), .ZN(n1290) );
  AO21X1 U1944 ( .IN1(n1803), .IN2(n1302), .IN3(n2046), .Q(n1466) );
  XOR2X1 U1945 ( .IN1(keyinput28), .IN2(n2047), .Q(n2046) );
  NOR2X0 U1946 ( .IN1(n1803), .IN2(n2048), .QN(n2047) );
  XNOR2X1 U1947 ( .IN1(keyinput11), .IN2(n1302), .Q(n2048) );
  INVX0 U1948 ( .INP(n1303), .ZN(n1803) );
  NAND3X0 U1949 ( .IN1(n1457), .IN2(n2049), .IN3(n2050), .QN(n1467) );
  OR4X1 U1950 ( .IN1(n1455), .IN2(n1445), .IN3(n1452), .IN4(n1434), .Q(n2050)
         );
  INVX0 U1951 ( .INP(n1437), .ZN(n1434) );
  AO21X1 U1952 ( .IN1(n1359), .IN2(n2051), .IN3(n1512), .Q(n1437) );
  NAND2X0 U1953 ( .IN1(n1490), .IN2(n2052), .QN(n2051) );
  NAND3X0 U1954 ( .IN1(n2053), .IN2(n1477), .IN3(n1352), .QN(n2052) );
  AO22X1 U1955 ( .IN1(n1544), .IN2(n2054), .IN3(n2055), .IN4(n1541), .Q(n1477)
         );
  NOR2X0 U1956 ( .IN1(keyinput31), .IN2(n1379), .QN(n2055) );
  OR2X1 U1957 ( .IN1(n1394), .IN2(keyinput31), .Q(n2054) );
  NAND2X0 U1958 ( .IN1(n1376), .IN2(n1495), .QN(n2053) );
  INVX0 U1959 ( .INP(n1479), .ZN(n1495) );
  NOR2X0 U1960 ( .IN1(n1370), .IN2(n1485), .QN(n1479) );
  AOI22X1 U1961 ( .IN1(n1515), .IN2(n1516), .IN3(n1237), .IN4(n2056), .QN(
        n1485) );
  NAND2X0 U1962 ( .IN1(n2057), .IN2(n2058), .QN(n2056) );
  NAND3X0 U1963 ( .IN1(n1268), .IN2(n2059), .IN3(n1403), .QN(n2058) );
  AO21X1 U1964 ( .IN1(n1412), .IN2(n2060), .IN3(n1414), .Q(n2059) );
  NOR2X0 U1965 ( .IN1(n1537), .IN2(N352), .QN(n1414) );
  INVX0 U1966 ( .INP(n2061), .ZN(n1537) );
  AO21X1 U1967 ( .IN1(n1225), .IN2(n2062), .IN3(n1425), .Q(n2060) );
  NAND4X0 U1968 ( .IN1(n2063), .IN2(n1227), .IN3(n1228), .IN4(n1229), .QN(
        n1425) );
  NAND3X0 U1969 ( .IN1(n1539), .IN2(n1419), .IN3(n1205), .QN(n1228) );
  INVX0 U1970 ( .INP(n1208), .ZN(n1539) );
  NAND2X0 U1971 ( .IN1(n1207), .IN2(n1419), .QN(n1227) );
  INVX0 U1972 ( .INP(n1210), .ZN(n1207) );
  NAND2X0 U1973 ( .IN1(n1230), .IN2(n2064), .QN(n2063) );
  NAND3X0 U1974 ( .IN1(n1426), .IN2(n1427), .IN3(n2065), .QN(n2062) );
  NAND2X0 U1975 ( .IN1(n1272), .IN2(n1430), .QN(n2065) );
  AO221X1 U1976 ( .IN1(n1141), .IN2(n2066), .IN3(n1526), .IN4(n1854), .IN5(
        n1527), .Q(n1430) );
  AND2X1 U1977 ( .IN1(n1856), .IN2(n1141), .Q(n1526) );
  NOR2X0 U1978 ( .IN1(n1128), .IN2(n1149), .QN(n1856) );
  OR2X1 U1979 ( .IN1(n1155), .IN2(n1529), .Q(n1149) );
  OR2X1 U1980 ( .IN1(n1131), .IN2(n1159), .Q(n1155) );
  INVX0 U1981 ( .INP(N367), .ZN(n1128) );
  AO21X1 U1982 ( .IN1(n1857), .IN2(n1854), .IN3(n1861), .Q(n2066) );
  NOR2X0 U1983 ( .IN1(n1533), .IN2(N319), .QN(n1861) );
  INVX0 U1984 ( .INP(n2067), .ZN(n1533) );
  AO21X1 U1985 ( .IN1(N319), .IN2(n2067), .IN3(n2068), .Q(n1854) );
  XOR2X1 U1986 ( .IN1(n2069), .IN2(keyinput63), .Q(n2068) );
  OR2X1 U1987 ( .IN1(n2067), .IN2(N319), .Q(n2069) );
  MUX21X1 U1988 ( .IN1(N236), .IN2(N23), .S(n1122), .Q(n2067) );
  AO21X1 U1989 ( .IN1(n1158), .IN2(n2070), .IN3(n1862), .Q(n1857) );
  OAI21X1 U1990 ( .IN1(n1138), .IN2(n1159), .IN3(n1863), .QN(n2070) );
  XNOR2X1 U1991 ( .IN1(n1532), .IN2(keyinput34), .Q(n1863) );
  AO21X1 U1992 ( .IN1(N313), .IN2(n1818), .IN3(n1532), .Q(n1159) );
  NOR2X0 U1993 ( .IN1(n1818), .IN2(N313), .QN(n1532) );
  INVX0 U1994 ( .INP(n2071), .ZN(n1818) );
  MUX21X1 U1995 ( .IN1(N238), .IN2(N29), .S(n1121), .Q(n2071) );
  INVX0 U1996 ( .INP(n1529), .ZN(n1158) );
  AO21X1 U1997 ( .IN1(n2072), .IN2(n1966), .IN3(n1862), .Q(n1529) );
  NOR2X0 U1998 ( .IN1(n1966), .IN2(n2072), .QN(n1862) );
  XOR2X1 U1999 ( .IN1(keyinput3), .IN2(N316), .Q(n1966) );
  INVX0 U2000 ( .INP(n1819), .ZN(n2072) );
  MUX21X1 U2001 ( .IN1(N237), .IN2(N26), .S(n1120), .Q(n1819) );
  INVX0 U2002 ( .INP(n1156), .ZN(n1141) );
  AO21X1 U2003 ( .IN1(N322), .IN2(n2073), .IN3(n1527), .Q(n1156) );
  NOR2X0 U2004 ( .IN1(n2073), .IN2(N322), .QN(n1527) );
  INVX0 U2005 ( .INP(n1812), .ZN(n2073) );
  MUX21X1 U2006 ( .IN1(N235), .IN2(N103), .S(n1119), .Q(n1812) );
  AND3X1 U2007 ( .IN1(n1184), .IN2(n1174), .IN3(n1175), .Q(n1272) );
  NOR2X0 U2008 ( .IN1(n1834), .IN2(n1183), .QN(n1175) );
  INVX0 U2009 ( .INP(n1172), .ZN(n1834) );
  NOR2X0 U2010 ( .IN1(n1182), .IN2(n1179), .QN(n1172) );
  NOR2X0 U2011 ( .IN1(n1984), .IN2(n1811), .QN(n1179) );
  INVX0 U2012 ( .INP(n1161), .ZN(n1174) );
  INVX0 U2013 ( .INP(n1850), .ZN(n1426) );
  OA21X1 U2014 ( .IN1(n1844), .IN2(n1522), .IN3(n1184), .Q(n1850) );
  OA21X1 U2015 ( .IN1(n1981), .IN2(n1805), .IN3(n1427), .Q(n1184) );
  NAND2X0 U2016 ( .IN1(n1805), .IN2(n1981), .QN(n1427) );
  MUX21X1 U2017 ( .IN1(N231), .IN2(N100), .S(n1122), .Q(n1805) );
  INVX0 U2018 ( .INP(N334), .ZN(n1981) );
  NOR2X0 U2019 ( .IN1(n1161), .IN2(n1843), .QN(n1844) );
  OA21X1 U2020 ( .IN1(n1183), .IN2(n1837), .IN3(n2074), .Q(n1843) );
  XNOR2X1 U2021 ( .IN1(keyinput32), .IN2(n1524), .Q(n2074) );
  XNOR2X1 U2022 ( .IN1(n1182), .IN2(keyinput33), .Q(n1837) );
  AND2X1 U2023 ( .IN1(n1811), .IN2(n1984), .Q(n1182) );
  XOR2X1 U2024 ( .IN1(keyinput4), .IN2(N325), .Q(n1984) );
  MUX21X1 U2025 ( .IN1(N234), .IN2(N130), .S(n1121), .Q(n1811) );
  AO21X1 U2026 ( .IN1(n1976), .IN2(n1809), .IN3(n1524), .Q(n1183) );
  NOR2X0 U2027 ( .IN1(n1809), .IN2(n1976), .QN(n1524) );
  INVX0 U2028 ( .INP(n2075), .ZN(n1809) );
  MUX21X1 U2029 ( .IN1(N233), .IN2(N127), .S(n1120), .Q(n2075) );
  XNOR2X1 U2030 ( .IN1(keyinput5), .IN2(N328), .Q(n1976) );
  AO21X1 U2031 ( .IN1(N331), .IN2(n1804), .IN3(n1522), .Q(n1161) );
  NOR2X0 U2032 ( .IN1(n1804), .IN2(N331), .QN(n1522) );
  INVX0 U2033 ( .INP(n2076), .ZN(n1804) );
  MUX21X1 U2034 ( .IN1(N232), .IN2(N124), .S(n1119), .Q(n2076) );
  AND2X1 U2035 ( .IN1(n1423), .IN2(n1230), .Q(n1225) );
  AND3X1 U2036 ( .IN1(n1205), .IN2(n1419), .IN3(n1224), .Q(n1230) );
  OA21X1 U2037 ( .IN1(n2005), .IN2(n1833), .IN3(n1208), .Q(n1224) );
  NAND2X0 U2038 ( .IN1(n1833), .IN2(n2005), .QN(n1208) );
  MUX21X1 U2039 ( .IN1(N226), .IN2(N97), .S(n1122), .Q(n1833) );
  INVX0 U2040 ( .INP(N343), .ZN(n2005) );
  OA21X1 U2041 ( .IN1(n2006), .IN2(n1830), .IN3(n1229), .Q(n1419) );
  NAND2X0 U2042 ( .IN1(n1830), .IN2(n2006), .QN(n1229) );
  MUX21X1 U2043 ( .IN1(N224), .IN2(N121), .S(n1121), .Q(n1830) );
  INVX0 U2044 ( .INP(N349), .ZN(n2006) );
  OA21X1 U2045 ( .IN1(n2004), .IN2(n1832), .IN3(n1210), .Q(n1205) );
  NAND2X0 U2046 ( .IN1(n1832), .IN2(n2004), .QN(n1210) );
  MUX21X1 U2047 ( .IN1(N225), .IN2(N94), .S(n1120), .Q(n1832) );
  INVX0 U2048 ( .INP(N346), .ZN(n2004) );
  NOR2X0 U2049 ( .IN1(n1222), .IN2(n2064), .QN(n1423) );
  INVX0 U2050 ( .INP(n1422), .ZN(n2064) );
  NAND2X0 U2051 ( .IN1(n1827), .IN2(n2002), .QN(n1422) );
  NOR2X0 U2052 ( .IN1(n2002), .IN2(n1827), .QN(n1222) );
  MUX21X1 U2053 ( .IN1(N217), .IN2(N118), .S(n1119), .Q(n1827) );
  INVX0 U2054 ( .INP(N340), .ZN(n2002) );
  XNOR2X1 U2055 ( .IN1(N352), .IN2(n2061), .Q(n1412) );
  MUX21X1 U2056 ( .IN1(N223), .IN2(N47), .S(n1122), .Q(n2061) );
  INVX0 U2057 ( .INP(n1264), .ZN(n1268) );
  NAND2X0 U2058 ( .IN1(n1249), .IN2(n1248), .QN(n1264) );
  NOR2X0 U2059 ( .IN1(n1251), .IN2(n2077), .QN(n1249) );
  INVX0 U2060 ( .INP(n1267), .ZN(n2077) );
  NAND2X0 U2061 ( .IN1(N355), .IN2(n1828), .QN(n1267) );
  INVX0 U2062 ( .INP(n1408), .ZN(n2057) );
  AO21X1 U2063 ( .IN1(n1403), .IN2(n1404), .IN3(n1540), .Q(n1408) );
  INVX0 U2064 ( .INP(n1242), .ZN(n1540) );
  NAND2X0 U2065 ( .IN1(n2078), .IN2(n1247), .QN(n1404) );
  NAND2X0 U2066 ( .IN1(n1251), .IN2(n1248), .QN(n1247) );
  OA21X1 U2067 ( .IN1(n1992), .IN2(n1829), .IN3(n1245), .Q(n1248) );
  NOR2X0 U2068 ( .IN1(n1828), .IN2(N355), .QN(n1251) );
  INVX0 U2069 ( .INP(n2079), .ZN(n1828) );
  MUX21X1 U2070 ( .IN1(N222), .IN2(N35), .S(n1121), .Q(n2079) );
  XOR2X1 U2071 ( .IN1(n1245), .IN2(keyinput37), .Q(n2078) );
  NAND2X0 U2072 ( .IN1(n1829), .IN2(n1992), .QN(n1245) );
  INVX0 U2073 ( .INP(N358), .ZN(n1992) );
  MUX21X1 U2074 ( .IN1(N221), .IN2(N32), .S(n1120), .Q(n1829) );
  MUX21X1 U2075 ( .IN1(n1252), .IN2(n2080), .S(keyinput58), .Q(n1403) );
  NAND2X0 U2076 ( .IN1(N361), .IN2(n1821), .QN(n2080) );
  OA21X1 U2077 ( .IN1(n1987), .IN2(n1821), .IN3(n1242), .Q(n1252) );
  NAND2X0 U2078 ( .IN1(n1821), .IN2(n1987), .QN(n1242) );
  MUX21X1 U2079 ( .IN1(N220), .IN2(N50), .S(n1119), .Q(n1821) );
  INVX0 U2080 ( .INP(N361), .ZN(n1987) );
  XNOR2X1 U2081 ( .IN1(N364), .IN2(n1515), .Q(n1237) );
  INVX0 U2082 ( .INP(N364), .ZN(n1516) );
  MUX21X1 U2083 ( .IN1(N66), .IN2(N219), .S(N18), .Q(n1515) );
  INVX0 U2084 ( .INP(n1381), .ZN(n1370) );
  NOR2X0 U2085 ( .IN1(n1386), .IN2(n1369), .QN(n1381) );
  INVX0 U2086 ( .INP(n1367), .ZN(n1386) );
  OA21X1 U2087 ( .IN1(n1919), .IN2(n2081), .IN3(n1486), .Q(n1367) );
  INVX0 U2088 ( .INP(N277), .ZN(n1919) );
  INVX0 U2089 ( .INP(n1382), .ZN(n1376) );
  NAND2X0 U2090 ( .IN1(n1393), .IN2(n1389), .QN(n1382) );
  INVX0 U2091 ( .INP(n1493), .ZN(n1389) );
  NOR2X0 U2092 ( .IN1(n1486), .IN2(n1369), .QN(n1493) );
  INVX0 U2093 ( .INP(n1475), .ZN(n1369) );
  OA21X1 U2094 ( .IN1(n1913), .IN2(n1782), .IN3(n1393), .Q(n1475) );
  INVX0 U2095 ( .INP(n1391), .ZN(n1486) );
  NOR2X0 U2096 ( .IN1(n1384), .IN2(N277), .QN(n1391) );
  INVX0 U2097 ( .INP(n2081), .ZN(n1384) );
  MUX21X1 U2098 ( .IN1(N151), .IN2(N147), .S(n1122), .Q(n2081) );
  NAND2X0 U2099 ( .IN1(n1782), .IN2(n1913), .QN(n1393) );
  INVX0 U2100 ( .INP(N280), .ZN(n1913) );
  MUX21X1 U2101 ( .IN1(N160), .IN2(N138), .S(n1121), .Q(n1782) );
  AOI21X1 U2102 ( .IN1(n1352), .IN2(n1379), .IN3(n2082), .QN(n1490) );
  INVX0 U2103 ( .INP(n1394), .ZN(n1379) );
  NAND2X0 U2104 ( .IN1(n1541), .IN2(n1544), .QN(n1394) );
  MUX21X1 U2105 ( .IN1(N144), .IN2(N159), .S(N18), .Q(n1544) );
  XNOR2X1 U2106 ( .IN1(keyinput2), .IN2(N283), .Q(n1541) );
  AOI21X1 U2107 ( .IN1(N286), .IN2(n2083), .IN3(n2082), .QN(n1352) );
  NOR2X0 U2108 ( .IN1(n2083), .IN2(N286), .QN(n2082) );
  INVX0 U2109 ( .INP(n1788), .ZN(n2083) );
  MUX21X1 U2110 ( .IN1(N158), .IN2(N135), .S(n1120), .Q(n1788) );
  AOI21X1 U2111 ( .IN1(N289), .IN2(n1787), .IN3(n1512), .QN(n1359) );
  NOR2X0 U2112 ( .IN1(n1787), .IN2(N289), .QN(n1512) );
  AOI21X1 U2113 ( .IN1(N157), .IN2(n1801), .IN3(n1802), .QN(n1787) );
  NAND2X0 U2114 ( .IN1(n1435), .IN2(n1442), .QN(n1455) );
  AND2X1 U2115 ( .IN1(n1339), .IN2(n1348), .Q(n1435) );
  INVX0 U2116 ( .INP(n1443), .ZN(n1348) );
  NAND2X0 U2117 ( .IN1(N293), .IN2(n1773), .QN(n1339) );
  INVX0 U2118 ( .INP(n1509), .ZN(n2049) );
  NAND2X0 U2119 ( .IN1(n1323), .IN2(n1456), .QN(n1457) );
  AO21X1 U2120 ( .IN1(n1453), .IN2(n2084), .IN3(n1454), .Q(n1456) );
  NAND2X0 U2121 ( .IN1(n1441), .IN2(n1446), .QN(n2084) );
  OR2X1 U2122 ( .IN1(N296), .IN2(n1546), .Q(n1446) );
  NAND2X0 U2123 ( .IN1(n1443), .IN2(n1442), .QN(n1441) );
  XNOR2X1 U2124 ( .IN1(n1546), .IN2(n1920), .Q(n1442) );
  INVX0 U2125 ( .INP(N296), .ZN(n1920) );
  AOI21X1 U2126 ( .IN1(N155), .IN2(n1801), .IN3(n1802), .QN(n1546) );
  NOR2X0 U2127 ( .IN1(n1773), .IN2(N293), .QN(n1443) );
  AOI21X1 U2128 ( .IN1(N156), .IN2(n1801), .IN3(n1802), .QN(n1773) );
  INVX0 U2129 ( .INP(n1445), .ZN(n1453) );
  AO21X1 U2130 ( .IN1(N299), .IN2(n2085), .IN3(n1454), .Q(n1445) );
  NOR2X0 U2131 ( .IN1(N299), .IN2(n2085), .QN(n1454) );
  INVX0 U2132 ( .INP(n1548), .ZN(n2085) );
  AO21X1 U2133 ( .IN1(N154), .IN2(n1801), .IN3(n1802), .Q(n1548) );
  INVX0 U2134 ( .INP(n1452), .ZN(n1323) );
  AO21X1 U2135 ( .IN1(N303), .IN2(n1791), .IN3(n1509), .Q(n1452) );
  NOR2X0 U2136 ( .IN1(n1791), .IN2(N303), .QN(n1509) );
  AOI21X1 U2137 ( .IN1(N153), .IN2(n1801), .IN3(n1802), .QN(n1791) );
  OA21X1 U2138 ( .IN1(n1296), .IN2(n1288), .IN3(n2086), .Q(n1294) );
  INVX0 U2139 ( .INP(n1291), .ZN(n2086) );
  NAND2X0 U2140 ( .IN1(n1302), .IN2(n1303), .QN(n1288) );
  AO21X1 U2141 ( .IN1(N209), .IN2(n1801), .IN3(n1802), .Q(n1303) );
  INVX0 U2142 ( .INP(N251), .ZN(n1302) );
  AO21X1 U2143 ( .IN1(N254), .IN2(n1794), .IN3(n1291), .Q(n1296) );
  NOR2X0 U2144 ( .IN1(N254), .IN2(n1794), .QN(n1291) );
  AOI21X1 U2145 ( .IN1(N216), .IN2(n1801), .IN3(n1802), .QN(n1794) );
  XNOR2X1 U2146 ( .IN1(n1503), .IN2(N106), .Q(n1469) );
  OA21X1 U2147 ( .IN1(n1306), .IN2(n1474), .IN3(n1473), .Q(n1311) );
  INVX0 U2148 ( .INP(n2087), .ZN(n1473) );
  NAND2X0 U2149 ( .IN1(n2032), .IN2(n1503), .QN(n1474) );
  AO21X1 U2150 ( .IN1(N215), .IN2(n1801), .IN3(n1802), .Q(n1503) );
  INVX0 U2151 ( .INP(N106), .ZN(n2032) );
  AO21X1 U2152 ( .IN1(N257), .IN2(n1797), .IN3(n2087), .Q(n1306) );
  NOR2X0 U2153 ( .IN1(N257), .IN2(n1797), .QN(n2087) );
  AOI21X1 U2154 ( .IN1(N214), .IN2(n1801), .IN3(n1802), .QN(n1797) );
  AND2X1 U2155 ( .IN1(n1801), .IN2(n1120), .Q(n1802) );
  XNOR2X1 U2156 ( .IN1(n1588), .IN2(keyinput1), .Q(n1801) );
  NAND2X0 U2157 ( .IN1(N9), .IN2(N12), .QN(n1588) );
  NOR2X0 U2158 ( .IN1(n1319), .IN2(n1318), .QN(n1320) );
  XOR2X1 U2159 ( .IN1(n2041), .IN2(n2018), .Q(n1318) );
  NAND2X0 U2160 ( .IN1(N267), .IN2(N382), .QN(n2041) );
  NAND2X0 U2161 ( .IN1(n1317), .IN2(n1316), .QN(n1319) );
  NAND3X0 U2162 ( .IN1(N263), .IN2(n2018), .IN3(N382), .QN(n1316) );
  AO21X1 U2163 ( .IN1(N382), .IN2(N263), .IN3(n2018), .Q(n1317) );
  INVX0 U2164 ( .INP(N38), .ZN(n2018) );
  XNOR2X1 U2165 ( .IN1(N367), .IN2(n1131), .Q(N10025) );
  NAND2X0 U2166 ( .IN1(n1154), .IN2(n1138), .QN(n1131) );
  NAND3X0 U2167 ( .IN1(n2088), .IN2(n1122), .IN3(n1817), .QN(n1138) );
  AO21X1 U2168 ( .IN1(n1817), .IN2(n1121), .IN3(n2088), .Q(n1154) );
  XNOR2X1 U2169 ( .IN1(n2089), .IN2(keyinput19), .Q(n2088) );
  NAND2X0 U2170 ( .IN1(N310), .IN2(n1119), .QN(n2089) );
  MUX21X1 U2171 ( .IN1(N229), .IN2(N41), .S(n1119), .Q(n1817) );
endmodule

