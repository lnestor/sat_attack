
module c2670 ( N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, 
        N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, 
        N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, 
        N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, 
        N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, 
        N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, 
        N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, 
        N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, 
        N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, 
        N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, 
        N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, 
        N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, 
        N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I, N149_I, 
        N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, 
        N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, 
        N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, 
        N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I, 
        N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, 
        N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, 
        N204_I, N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, 
        N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, N401, N419, 
        N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, 
        N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, 
        N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, 
        N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, 
        N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, 
        N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, N144_O, 
        N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, 
        N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, 
        N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, 
        N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, 
        N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, 
        N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, 
        N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O, 
        N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, 
        N217_O, N218_O, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31 );
  input N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40,
         N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227,
         N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263,
         N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297,
         N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334,
         N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I,
         N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I,
         N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I,
         N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I,
         N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, N177_I,
         N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I,
         N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I,
         N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I,
         N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I,
         N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, N217_I,
         N218_I, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
         keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10,
         keyinput11, keyinput12, keyinput13, keyinput14, keyinput15,
         keyinput16, keyinput17, keyinput18, keyinput19, keyinput20,
         keyinput21, keyinput22, keyinput23, keyinput24, keyinput25,
         keyinput26, keyinput27, keyinput28, keyinput29, keyinput30,
         keyinput31;
  output N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489,
         N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029,
         N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821,
         N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022,
         N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970,
         N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875,
         N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O,
         N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O,
         N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O,
         N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O,
         N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O,
         N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O,
         N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O,
         N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O,
         N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O,
         N214_O, N215_O, N216_O, N217_O, N218_O;
  wire   N219, N253, N290, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I,
         N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I,
         N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I,
         N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I,
         N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I,
         N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I,
         N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I,
         N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I,
         N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I,
         N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N2387, N2389, N2643,
         N3803, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600;
  assign N805 = N219;
  assign N401 = N219;
  assign N400 = N219;
  assign N398 = N219;
  assign N420 = N253;
  assign N419 = N253;
  assign N458 = N290;
  assign N457 = N290;
  assign N456 = N290;
  assign N143_O = N143_I;
  assign N144_O = N144_I;
  assign N145_O = N145_I;
  assign N146_O = N146_I;
  assign N147_O = N147_I;
  assign N148_O = N148_I;
  assign N149_O = N149_I;
  assign N150_O = N150_I;
  assign N151_O = N151_I;
  assign N152_O = N152_I;
  assign N153_O = N153_I;
  assign N154_O = N154_I;
  assign N155_O = N155_I;
  assign N156_O = N156_I;
  assign N157_O = N157_I;
  assign N158_O = N158_I;
  assign N159_O = N159_I;
  assign N160_O = N160_I;
  assign N161_O = N161_I;
  assign N162_O = N162_I;
  assign N163_O = N163_I;
  assign N164_O = N164_I;
  assign N165_O = N165_I;
  assign N166_O = N166_I;
  assign N167_O = N167_I;
  assign N168_O = N168_I;
  assign N169_O = N169_I;
  assign N170_O = N170_I;
  assign N171_O = N171_I;
  assign N172_O = N172_I;
  assign N173_O = N173_I;
  assign N174_O = N174_I;
  assign N175_O = N175_I;
  assign N176_O = N176_I;
  assign N177_O = N177_I;
  assign N178_O = N178_I;
  assign N179_O = N179_I;
  assign N180_O = N180_I;
  assign N181_O = N181_I;
  assign N182_O = N182_I;
  assign N183_O = N183_I;
  assign N184_O = N184_I;
  assign N185_O = N185_I;
  assign N186_O = N186_I;
  assign N187_O = N187_I;
  assign N188_O = N188_I;
  assign N189_O = N189_I;
  assign N190_O = N190_I;
  assign N191_O = N191_I;
  assign N192_O = N192_I;
  assign N193_O = N193_I;
  assign N194_O = N194_I;
  assign N195_O = N195_I;
  assign N196_O = N196_I;
  assign N197_O = N197_I;
  assign N198_O = N198_I;
  assign N199_O = N199_I;
  assign N200_O = N200_I;
  assign N201_O = N201_I;
  assign N202_O = N202_I;
  assign N203_O = N203_I;
  assign N204_O = N204_I;
  assign N205_O = N205_I;
  assign N206_O = N206_I;
  assign N207_O = N207_I;
  assign N208_O = N208_I;
  assign N209_O = N209_I;
  assign N210_O = N210_I;
  assign N211_O = N211_I;
  assign N212_O = N212_I;
  assign N213_O = N213_I;
  assign N214_O = N214_I;
  assign N215_O = N215_I;
  assign N216_O = N216_I;
  assign N217_O = N217_I;
  assign N218_O = N218_I;
  assign N2388 = N2387;
  assign N2390 = N2389;
  assign N2644 = N2643;
  assign N3804 = N3803;

  NAND3X0 U364 ( .IN1(N2), .IN2(N15), .IN3(N237), .QN(N799) );
  NAND4X0 U365 ( .IN1(N309), .IN2(N305), .IN3(N301), .IN4(N297), .QN(N792) );
  INVX0 U366 ( .INP(N108), .ZN(N494) );
  INVX0 U367 ( .INP(N57), .ZN(N493) );
  INVX0 U368 ( .INP(N120), .ZN(N492) );
  INVX0 U369 ( .INP(N69), .ZN(N491) );
  INVX0 U370 ( .INP(N96), .ZN(N490) );
  INVX0 U371 ( .INP(N82), .ZN(N489) );
  INVX0 U372 ( .INP(N132), .ZN(N488) );
  INVX0 U373 ( .INP(N44), .ZN(N487) );
  INVX0 U374 ( .INP(N3882), .ZN(N3881) );
  NAND4X0 U375 ( .IN1(n340), .IN2(n341), .IN3(N1726), .IN4(n342), .QN(N3882)
         );
  NOR4X0 U376 ( .IN1(N3809), .IN2(N3671), .IN3(N2925), .IN4(N2970), .QN(n342)
         );
  INVX0 U377 ( .INP(N3875), .ZN(n340) );
  XNOR2X1 U378 ( .IN1(N3851), .IN2(n343), .Q(N3875) );
  OA21X1 U379 ( .IN1(keyinput31), .IN2(n344), .IN3(n345), .Q(n343) );
  AO22X1 U380 ( .IN1(n344), .IN2(n346), .IN3(n347), .IN4(n348), .Q(n345) );
  OR4X1 U381 ( .IN1(n349), .IN2(n350), .IN3(n351), .IN4(n352), .Q(n348) );
  OR3X1 U382 ( .IN1(n353), .IN2(n354), .IN3(n355), .Q(n352) );
  OA22X1 U383 ( .IN1(n356), .IN2(n357), .IN3(N2010), .IN4(n358), .Q(n354) );
  NOR2X0 U384 ( .IN1(n359), .IN2(n360), .QN(n356) );
  XOR2X1 U385 ( .IN1(n361), .IN2(keyinput24), .Q(n360) );
  XOR2X1 U386 ( .IN1(keyinput30), .IN2(n362), .Q(n347) );
  OA21X1 U387 ( .IN1(n363), .IN2(n349), .IN3(n364), .Q(n362) );
  OA21X1 U388 ( .IN1(n365), .IN2(n350), .IN3(n366), .Q(n363) );
  OA21X1 U389 ( .IN1(n367), .IN2(n353), .IN3(n368), .Q(n365) );
  OA22X1 U390 ( .IN1(n351), .IN2(n369), .IN3(n370), .IN4(n371), .Q(n367) );
  XNOR2X1 U391 ( .IN1(n370), .IN2(n371), .Q(n351) );
  OR2X1 U392 ( .IN1(n372), .IN2(n373), .Q(n371) );
  NAND4X0 U393 ( .IN1(n374), .IN2(n375), .IN3(n376), .IN4(n377), .QN(n346) );
  NAND2X0 U394 ( .IN1(n378), .IN2(n379), .QN(n374) );
  AOI21X1 U395 ( .IN1(n380), .IN2(n377), .IN3(n381), .QN(n344) );
  AO22X1 U396 ( .IN1(n382), .IN2(n383), .IN3(n376), .IN4(n384), .Q(n380) );
  NAND2X0 U397 ( .IN1(n385), .IN2(n386), .QN(n384) );
  INVX0 U398 ( .INP(n387), .ZN(n386) );
  NAND3X0 U399 ( .IN1(n388), .IN2(n375), .IN3(n389), .QN(n385) );
  INVX0 U400 ( .INP(n379), .ZN(n389) );
  NAND2X0 U401 ( .IN1(n390), .IN2(n391), .QN(n379) );
  XNOR2X1 U402 ( .IN1(N281), .IN2(keyinput21), .Q(n390) );
  OR2X1 U403 ( .IN1(n383), .IN2(n382), .Q(n376) );
  AO21X1 U404 ( .IN1(n392), .IN2(n393), .IN3(n381), .Q(N3851) );
  NOR3X0 U405 ( .IN1(n394), .IN2(N294), .IN3(n395), .QN(n381) );
  AO22X1 U406 ( .IN1(n382), .IN2(n396), .IN3(n397), .IN4(n398), .Q(n393) );
  NOR2X0 U407 ( .IN1(keyinput27), .IN2(n399), .QN(n397) );
  NAND2X0 U408 ( .IN1(n399), .IN2(n400), .QN(n396) );
  INVX0 U409 ( .INP(n398), .ZN(n400) );
  XNOR2X1 U410 ( .IN1(n383), .IN2(keyinput20), .Q(n398) );
  NAND2X0 U411 ( .IN1(n391), .IN2(n401), .QN(n383) );
  AOI21X1 U412 ( .IN1(n402), .IN2(n375), .IN3(n387), .QN(n399) );
  NOR3X0 U413 ( .IN1(n403), .IN2(N284), .IN3(n395), .QN(n387) );
  NAND3X0 U414 ( .IN1(N284), .IN2(n403), .IN3(n391), .QN(n375) );
  AO22X1 U415 ( .IN1(n388), .IN2(n404), .IN3(n405), .IN4(n391), .Q(n402) );
  NOR2X0 U416 ( .IN1(N281), .IN2(n406), .QN(n405) );
  OA21X1 U417 ( .IN1(keyinput26), .IN2(n407), .IN3(n378), .Q(n406) );
  INVX0 U418 ( .INP(n388), .ZN(n378) );
  INVX0 U419 ( .INP(n407), .ZN(n404) );
  OA21X1 U420 ( .IN1(n408), .IN2(n409), .IN3(n364), .Q(n407) );
  XNOR2X1 U421 ( .IN1(keyinput29), .IN2(n349), .Q(n409) );
  NAND2X0 U422 ( .IN1(n364), .IN2(n410), .QN(n349) );
  NAND3X0 U423 ( .IN1(N278), .IN2(N2020), .IN3(n411), .QN(n410) );
  NAND3X0 U424 ( .IN1(n412), .IN2(n413), .IN3(n411), .QN(n364) );
  OA21X1 U425 ( .IN1(n414), .IN2(n350), .IN3(n366), .Q(n408) );
  NAND2X0 U426 ( .IN1(n366), .IN2(n415), .QN(n350) );
  NAND3X0 U427 ( .IN1(N275), .IN2(N2018), .IN3(n411), .QN(n415) );
  NAND3X0 U428 ( .IN1(n416), .IN2(n417), .IN3(n411), .QN(n366) );
  OA21X1 U429 ( .IN1(n418), .IN2(n353), .IN3(n368), .Q(n414) );
  NAND2X0 U430 ( .IN1(n368), .IN2(n419), .QN(n353) );
  OR3X1 U431 ( .IN1(n372), .IN2(N1819), .IN3(n420), .Q(n419) );
  NAND2X0 U432 ( .IN1(n420), .IN2(N1819), .QN(n368) );
  AO22X1 U433 ( .IN1(n411), .IN2(n421), .IN3(n422), .IN4(n423), .Q(n420) );
  NOR2X0 U434 ( .IN1(N309), .IN2(n372), .QN(n422) );
  INVX0 U435 ( .INP(N272), .ZN(n421) );
  NOR2X0 U436 ( .IN1(n372), .IN2(n423), .QN(n411) );
  OA22X1 U437 ( .IN1(n370), .IN2(n424), .IN3(n425), .IN4(n426), .Q(n418) );
  AND2X1 U438 ( .IN1(n424), .IN2(n370), .Q(n426) );
  OA21X1 U439 ( .IN1(n427), .IN2(n355), .IN3(n369), .Q(n425) );
  INVX0 U440 ( .INP(n428), .ZN(n369) );
  AO21X1 U441 ( .IN1(n429), .IN2(N2012), .IN3(n428), .Q(n355) );
  NOR2X0 U442 ( .IN1(n429), .IN2(N2012), .QN(n428) );
  MUX21X1 U443 ( .IN1(N301), .IN2(N266), .S(n430), .Q(n429) );
  OA22X1 U444 ( .IN1(n357), .IN2(n431), .IN3(N2010), .IN4(n358), .Q(n427) );
  AO22X1 U445 ( .IN1(n432), .IN2(N2010), .IN3(n433), .IN4(n361), .Q(n431) );
  MUX21X1 U446 ( .IN1(N287), .IN2(N256), .S(n430), .Q(n361) );
  INVX0 U447 ( .INP(keyinput14), .ZN(n432) );
  AO22X1 U448 ( .IN1(n358), .IN2(N2010), .IN3(n434), .IN4(n433), .Q(n357) );
  INVX0 U449 ( .INP(n359), .ZN(n433) );
  NOR2X0 U450 ( .IN1(n435), .IN2(n436), .QN(n359) );
  AO21X1 U451 ( .IN1(n435), .IN2(n436), .IN3(n437), .Q(n434) );
  MUX21X1 U452 ( .IN1(N294), .IN2(N259), .S(n430), .Q(n435) );
  MUX21X1 U453 ( .IN1(N263), .IN2(N297), .S(n423), .Q(n358) );
  INVX0 U454 ( .INP(n430), .ZN(n423) );
  NAND2X0 U455 ( .IN1(N8), .IN2(n438), .QN(n424) );
  XNOR2X1 U456 ( .IN1(keyinput25), .IN2(n373), .Q(n438) );
  MUX21X1 U457 ( .IN1(N305), .IN2(N269), .S(n430), .Q(n373) );
  NAND4X0 U458 ( .IN1(N40), .IN2(N1816), .IN3(n439), .IN4(n440), .QN(n430) );
  NOR2X0 U459 ( .IN1(n372), .IN2(N1820), .QN(n370) );
  INVX0 U460 ( .INP(N8), .ZN(n372) );
  NAND2X0 U461 ( .IN1(n391), .IN2(N2022), .QN(n388) );
  NOR2X0 U462 ( .IN1(n395), .IN2(N287), .QN(n382) );
  MUX21X1 U463 ( .IN1(n394), .IN2(n377), .S(keyinput28), .Q(n392) );
  NAND2X0 U464 ( .IN1(n394), .IN2(N294), .QN(n377) );
  AND2X1 U465 ( .IN1(n391), .IN2(n441), .Q(n394) );
  INVX0 U466 ( .INP(n395), .ZN(n391) );
  NAND3X0 U467 ( .IN1(N1816), .IN2(n442), .IN3(N40), .QN(n395) );
  NAND2X0 U468 ( .IN1(n439), .IN2(n440), .QN(n442) );
  INVX0 U469 ( .INP(N262), .ZN(n440) );
  AND2X1 U470 ( .IN1(n443), .IN2(n444), .Q(N3809) );
  XOR3X1 U471 ( .IN1(n445), .IN2(n446), .IN3(n447), .Q(n443) );
  NAND2X0 U472 ( .IN1(n448), .IN2(n449), .QN(n446) );
  XOR2X1 U473 ( .IN1(n450), .IN2(keyinput23), .Q(n449) );
  NAND3X0 U474 ( .IN1(n451), .IN2(n452), .IN3(n453), .QN(n450) );
  MUX21X1 U475 ( .IN1(n454), .IN2(n455), .S(n451), .Q(n448) );
  OR2X1 U476 ( .IN1(n452), .IN2(n453), .Q(n455) );
  XNOR2X1 U477 ( .IN1(n453), .IN2(n452), .Q(n454) );
  XNOR2X1 U478 ( .IN1(N1821), .IN2(N2014), .Q(n452) );
  AOI21X1 U479 ( .IN1(n436), .IN2(n456), .IN3(n457), .QN(n453) );
  XOR2X1 U480 ( .IN1(keyinput18), .IN2(n458), .Q(n457) );
  NOR2X0 U481 ( .IN1(n456), .IN2(n436), .QN(n458) );
  NOR2X0 U482 ( .IN1(keyinput22), .IN2(n459), .QN(n445) );
  MUX21X1 U483 ( .IN1(n460), .IN2(n461), .S(N246), .Q(N3803) );
  XOR2X1 U484 ( .IN1(n462), .IN2(n463), .Q(n461) );
  XNOR3X1 U485 ( .IN1(n464), .IN2(n456), .IN3(n436), .Q(n463) );
  XOR3X1 U486 ( .IN1(n451), .IN2(n459), .IN3(n447), .Q(n462) );
  XNOR2X1 U487 ( .IN1(N1819), .IN2(n416), .Q(n447) );
  XNOR2X1 U488 ( .IN1(N2022), .IN2(N2020), .Q(n459) );
  XNOR2X1 U489 ( .IN1(n437), .IN2(n460), .Q(n451) );
  AND2X1 U490 ( .IN1(n465), .IN2(n444), .Q(N3671) );
  INVX0 U491 ( .INP(N37), .ZN(n444) );
  XNOR3X1 U492 ( .IN1(n466), .IN2(n467), .IN3(n468), .Q(n465) );
  XNOR3X1 U493 ( .IN1(n469), .IN2(N1817), .IN3(n470), .Q(n468) );
  XNOR2X1 U494 ( .IN1(n471), .IN2(n472), .Q(n470) );
  AO221X1 U495 ( .IN1(N118), .IN2(n473), .IN3(N130), .IN4(n474), .IN5(n475), 
        .Q(n471) );
  AO22X1 U496 ( .IN1(N142), .IN2(n476), .IN3(N106), .IN4(n477), .Q(n475) );
  XNOR3X1 U497 ( .IN1(n401), .IN2(n441), .IN3(n478), .Q(n466) );
  XNOR2X1 U498 ( .IN1(n403), .IN2(n439), .Q(n478) );
  XNOR2X1 U499 ( .IN1(n479), .IN2(n460), .Q(N3546) );
  AO221X1 U500 ( .IN1(N67), .IN2(n480), .IN3(N55), .IN4(n481), .IN5(n482), .Q(
        n460) );
  AO22X1 U501 ( .IN1(N93), .IN2(n483), .IN3(N80), .IN4(n484), .Q(n482) );
  NAND2X0 U502 ( .IN1(n485), .IN2(n486), .QN(n479) );
  XNOR2X1 U503 ( .IN1(n437), .IN2(n487), .Q(n485) );
  NOR2X0 U504 ( .IN1(n464), .IN2(n436), .QN(n487) );
  XNOR2X1 U505 ( .IN1(n488), .IN2(n489), .Q(N2970) );
  XOR3X1 U506 ( .IN1(N305), .IN2(N294), .IN3(n490), .Q(n489) );
  OA21X1 U507 ( .IN1(N301), .IN2(n491), .IN3(n492), .Q(n490) );
  XOR2X1 U508 ( .IN1(n493), .IN2(keyinput2), .Q(n492) );
  NAND2X0 U509 ( .IN1(N301), .IN2(n491), .QN(n493) );
  XOR3X1 U510 ( .IN1(N313), .IN2(N309), .IN3(n494), .Q(n488) );
  XNOR2X1 U511 ( .IN1(N316), .IN2(N355), .Q(n494) );
  INVX0 U512 ( .INP(N3038), .ZN(N3079) );
  INVX0 U513 ( .INP(n341), .ZN(N2971) );
  XNOR3X1 U514 ( .IN1(N287), .IN2(N284), .IN3(n495), .Q(n341) );
  XOR3X1 U515 ( .IN1(n496), .IN2(n497), .IN3(n498), .Q(n495) );
  XNOR2X1 U516 ( .IN1(N263), .IN2(n499), .Q(n498) );
  OA21X1 U517 ( .IN1(N281), .IN2(n413), .IN3(n500), .Q(n499) );
  XOR2X1 U518 ( .IN1(keyinput3), .IN2(n501), .Q(n500) );
  AND2X1 U519 ( .IN1(n413), .IN2(N281), .Q(n501) );
  XNOR3X1 U520 ( .IN1(n417), .IN2(N272), .IN3(n502), .Q(n497) );
  XOR2X1 U521 ( .IN1(keyinput5), .IN2(N352), .Q(n502) );
  XOR2X1 U522 ( .IN1(N269), .IN2(N266), .Q(n496) );
  NOR4X0 U523 ( .IN1(n503), .IN2(n504), .IN3(n505), .IN4(n506), .QN(N3038) );
  NAND4X0 U524 ( .IN1(n507), .IN2(N11), .IN3(n508), .IN4(n509), .QN(n506) );
  XOR2X1 U525 ( .IN1(keyinput17), .IN2(n510), .Q(n509) );
  OA21X1 U526 ( .IN1(N301), .IN2(n511), .IN3(n512), .Q(n510) );
  XOR2X1 U527 ( .IN1(keyinput11), .IN2(n513), .Q(n512) );
  AND2X1 U528 ( .IN1(n511), .IN2(N301), .Q(n513) );
  MUX21X1 U529 ( .IN1(N27), .IN2(n439), .S(N29), .Q(n511) );
  XOR2X1 U530 ( .IN1(N309), .IN2(n514), .Q(n508) );
  MUX21X1 U531 ( .IN1(N35), .IN2(n515), .S(N29), .Q(n514) );
  XOR3X1 U532 ( .IN1(keyinput16), .IN2(N305), .IN3(n516), .Q(n507) );
  MUX21X1 U533 ( .IN1(N34), .IN2(n467), .S(N29), .Q(n516) );
  MUX21X1 U534 ( .IN1(n517), .IN2(n518), .S(N29), .Q(n505) );
  NAND2X0 U535 ( .IN1(n519), .IN2(n469), .QN(n518) );
  XOR2X1 U536 ( .IN1(n520), .IN2(n441), .Q(n519) );
  AO221X1 U537 ( .IN1(N116), .IN2(n473), .IN3(N128), .IN4(n474), .IN5(n521), 
        .Q(n441) );
  AO22X1 U538 ( .IN1(N140), .IN2(n476), .IN3(N104), .IN4(n477), .Q(n521) );
  NAND2X0 U539 ( .IN1(n522), .IN2(N28), .QN(n517) );
  XOR2X1 U540 ( .IN1(n520), .IN2(N26), .Q(n522) );
  OR2X1 U541 ( .IN1(keyinput10), .IN2(N294), .Q(n520) );
  MUX21X1 U542 ( .IN1(n523), .IN2(n524), .S(N29), .Q(n504) );
  NAND2X0 U543 ( .IN1(n525), .IN2(n526), .QN(n524) );
  XNOR2X1 U544 ( .IN1(n472), .IN2(n491), .Q(n526) );
  AO221X1 U545 ( .IN1(N139), .IN2(n476), .IN3(N115), .IN4(n473), .IN5(n527), 
        .Q(n472) );
  AO21X1 U546 ( .IN1(N127), .IN2(n474), .IN3(n528), .Q(n527) );
  XOR2X1 U547 ( .IN1(n529), .IN2(keyinput6), .Q(n528) );
  NAND2X0 U548 ( .IN1(N103), .IN2(n477), .QN(n529) );
  XOR2X1 U549 ( .IN1(n401), .IN2(N287), .Q(n525) );
  AO221X1 U550 ( .IN1(N117), .IN2(n473), .IN3(N129), .IN4(n474), .IN5(n530), 
        .Q(n401) );
  AO22X1 U551 ( .IN1(N141), .IN2(n476), .IN3(N105), .IN4(n477), .Q(n530) );
  NAND2X0 U552 ( .IN1(n531), .IN2(n532), .QN(n523) );
  XOR2X1 U553 ( .IN1(N32), .IN2(N287), .Q(n532) );
  XNOR2X1 U554 ( .IN1(N33), .IN2(n491), .Q(n531) );
  INVX0 U555 ( .INP(N297), .ZN(n491) );
  XNOR2X1 U556 ( .IN1(n533), .IN2(keyinput19), .Q(n503) );
  NAND3X0 U557 ( .IN1(n534), .IN2(n535), .IN3(n536), .QN(n533) );
  MUX21X1 U558 ( .IN1(n537), .IN2(n538), .S(N16), .Q(n536) );
  NOR2X0 U559 ( .IN1(n539), .IN2(n540), .QN(n538) );
  NAND4X0 U560 ( .IN1(n541), .IN2(n542), .IN3(n543), .IN4(n544), .QN(n540) );
  XNOR2X1 U561 ( .IN1(N1821), .IN2(N266), .Q(n544) );
  XNOR2X1 U562 ( .IN1(N1820), .IN2(N269), .Q(n543) );
  XNOR2X1 U563 ( .IN1(n416), .IN2(N275), .Q(n542) );
  INVX0 U564 ( .INP(N2018), .ZN(n416) );
  XNOR2X1 U565 ( .IN1(n412), .IN2(N278), .Q(n541) );
  INVX0 U566 ( .INP(N2020), .ZN(n412) );
  NAND4X0 U567 ( .IN1(n545), .IN2(n546), .IN3(n547), .IN4(n548), .QN(n539) );
  XOR2X1 U568 ( .IN1(n549), .IN2(N2022), .Q(n548) );
  XOR2X1 U569 ( .IN1(n436), .IN2(N259), .Q(n547) );
  XNOR2X1 U570 ( .IN1(n550), .IN2(N256), .Q(n546) );
  XNOR2X1 U571 ( .IN1(n456), .IN2(N263), .Q(n545) );
  INVX0 U572 ( .INP(N2010), .ZN(n456) );
  NOR2X0 U573 ( .IN1(n551), .IN2(n552), .QN(n537) );
  NAND4X0 U574 ( .IN1(n553), .IN2(n554), .IN3(n555), .IN4(n556), .QN(n552) );
  XOR2X1 U575 ( .IN1(N4), .IN2(N259), .Q(n556) );
  XOR2X1 U576 ( .IN1(N5), .IN2(N266), .Q(n555) );
  XNOR2X1 U577 ( .IN1(N6), .IN2(n413), .Q(n554) );
  INVX0 U578 ( .INP(N278), .ZN(n413) );
  XOR2X1 U579 ( .IN1(n549), .IN2(N24), .Q(n553) );
  OR2X1 U580 ( .IN1(keyinput9), .IN2(N281), .Q(n549) );
  NAND4X0 U581 ( .IN1(n557), .IN2(n558), .IN3(n559), .IN4(n560), .QN(n551) );
  XOR2X1 U582 ( .IN1(N256), .IN2(N19), .Q(n560) );
  XOR2X1 U583 ( .IN1(N263), .IN2(N20), .Q(n559) );
  XOR2X1 U584 ( .IN1(N269), .IN2(N21), .Q(n558) );
  XNOR2X1 U585 ( .IN1(n417), .IN2(N23), .Q(n557) );
  INVX0 U586 ( .INP(N275), .ZN(n417) );
  XNOR3X1 U587 ( .IN1(keyinput8), .IN2(n561), .IN3(N272), .Q(n535) );
  MUX21X1 U588 ( .IN1(N22), .IN2(N2016), .S(N16), .Q(n561) );
  XOR3X1 U589 ( .IN1(keyinput15), .IN2(N284), .IN3(n562), .Q(n534) );
  MUX21X1 U590 ( .IN1(N25), .IN2(n403), .S(N29), .Q(n562) );
  AO221X1 U591 ( .IN1(N107), .IN2(n473), .IN3(N119), .IN4(n474), .IN5(n563), 
        .Q(n403) );
  AO22X1 U592 ( .IN1(N131), .IN2(n476), .IN3(N95), .IN4(n477), .Q(n563) );
  NAND2X0 U593 ( .IN1(n564), .IN2(n565), .QN(N2891) );
  XNOR3X1 U594 ( .IN1(keyinput12), .IN2(N313), .IN3(n469), .Q(n565) );
  AO221X1 U595 ( .IN1(N111), .IN2(n473), .IN3(N123), .IN4(n474), .IN5(n566), 
        .Q(n469) );
  AO22X1 U596 ( .IN1(N135), .IN2(n476), .IN3(N99), .IN4(n477), .Q(n566) );
  XNOR2X1 U597 ( .IN1(N316), .IN2(keyinput7), .Q(n564) );
  AND2X1 U598 ( .IN1(N14), .IN2(n567), .Q(N2925) );
  XOR3X1 U599 ( .IN1(keyinput13), .IN2(N349), .IN3(n568), .Q(n567) );
  XOR3X1 U600 ( .IN1(n569), .IN2(n570), .IN3(N346), .Q(n568) );
  XOR3X1 U601 ( .IN1(N259), .IN2(N256), .IN3(n571), .Q(n570) );
  XOR2X1 U602 ( .IN1(N331), .IN2(N328), .Q(n571) );
  XOR3X1 U603 ( .IN1(N337), .IN2(N334), .IN3(n572), .Q(n569) );
  XOR2X1 U604 ( .IN1(N343), .IN2(N340), .Q(n572) );
  MUX21X1 U605 ( .IN1(n437), .IN2(n573), .S(N246), .Q(N2643) );
  AO21X1 U606 ( .IN1(n573), .IN2(n486), .IN3(n436), .Q(N2496) );
  INVX0 U607 ( .INP(N241), .ZN(n486) );
  INVX0 U608 ( .INP(n464), .ZN(n573) );
  NOR2X0 U609 ( .IN1(N230), .IN2(n436), .QN(n464) );
  MUX21X1 U610 ( .IN1(N2010), .IN2(N2014), .S(N246), .Q(N2389) );
  MUX21X1 U611 ( .IN1(n436), .IN2(N2012), .S(N246), .Q(N2387) );
  AO221X1 U612 ( .IN1(N66), .IN2(n480), .IN3(N54), .IN4(n481), .IN5(n574), .Q(
        n436) );
  AO22X1 U613 ( .IN1(N92), .IN2(n483), .IN3(N79), .IN4(n484), .Q(n574) );
  NAND2X0 U614 ( .IN1(n575), .IN2(n576), .QN(N1971) );
  XOR2X1 U615 ( .IN1(n577), .IN2(keyinput0), .Q(n575) );
  NAND2X0 U616 ( .IN1(N3), .IN2(N1), .QN(n577) );
  NAND2X0 U617 ( .IN1(N36), .IN2(n576), .QN(N1970) );
  AND3X1 U618 ( .IN1(N1726), .IN2(N237), .IN3(N224), .Q(n576) );
  NAND2X0 U619 ( .IN1(N241), .IN2(n550), .QN(N1969) );
  INVX0 U620 ( .INP(n437), .ZN(n550) );
  AO221X1 U621 ( .IN1(N56), .IN2(n480), .IN3(N43), .IN4(n481), .IN5(n578), .Q(
        n437) );
  AO22X1 U622 ( .IN1(N81), .IN2(n483), .IN3(N68), .IN4(n484), .Q(n578) );
  INVX0 U623 ( .INP(N2012), .ZN(N1821) );
  INVX0 U624 ( .INP(N2014), .ZN(N1820) );
  INVX0 U625 ( .INP(N2016), .ZN(N1819) );
  INVX0 U626 ( .INP(n439), .ZN(N1818) );
  AO221X1 U627 ( .IN1(N114), .IN2(n473), .IN3(N126), .IN4(n474), .IN5(n579), 
        .Q(n439) );
  AO22X1 U628 ( .IN1(N138), .IN2(n476), .IN3(N102), .IN4(n477), .Q(n579) );
  INVX0 U629 ( .INP(n515), .ZN(N1817) );
  AO221X1 U630 ( .IN1(N112), .IN2(n473), .IN3(N124), .IN4(n474), .IN5(n580), 
        .Q(n515) );
  AO22X1 U631 ( .IN1(N136), .IN2(n476), .IN3(N100), .IN4(n477), .Q(n580) );
  INVX0 U632 ( .INP(n467), .ZN(N1816) );
  AO221X1 U633 ( .IN1(N113), .IN2(n473), .IN3(N125), .IN4(n474), .IN5(n581), 
        .Q(n467) );
  AO22X1 U634 ( .IN1(N137), .IN2(n476), .IN3(N101), .IN4(n477), .Q(n581) );
  NOR2X0 U635 ( .IN1(n582), .IN2(N322), .QN(n477) );
  NOR2X0 U636 ( .IN1(N319), .IN2(N322), .QN(n476) );
  NOR2X0 U637 ( .IN1(n583), .IN2(N319), .QN(n474) );
  NOR2X0 U638 ( .IN1(n583), .IN2(n582), .QN(n473) );
  INVX0 U639 ( .INP(N319), .ZN(n582) );
  INVX0 U640 ( .INP(N322), .ZN(n583) );
  AO221X1 U641 ( .IN1(N60), .IN2(n480), .IN3(N47), .IN4(n481), .IN5(n584), .Q(
        N2022) );
  AO22X1 U642 ( .IN1(N85), .IN2(n483), .IN3(N72), .IN4(n484), .Q(n584) );
  AO221X1 U643 ( .IN1(N61), .IN2(n480), .IN3(N48), .IN4(n481), .IN5(n585), .Q(
        N2020) );
  AO22X1 U644 ( .IN1(N86), .IN2(n483), .IN3(N73), .IN4(n484), .Q(n585) );
  NAND4X0 U645 ( .IN1(n586), .IN2(n587), .IN3(n588), .IN4(n589), .QN(N2018) );
  NAND2X0 U646 ( .IN1(N87), .IN2(n590), .QN(n588) );
  NAND2X0 U647 ( .IN1(N74), .IN2(N234), .QN(n587) );
  XOR2X1 U648 ( .IN1(n591), .IN2(keyinput4), .Q(n586) );
  NAND2X0 U649 ( .IN1(N49), .IN2(n481), .QN(n591) );
  AO221X1 U650 ( .IN1(N88), .IN2(n483), .IN3(N62), .IN4(n480), .IN5(n592), .Q(
        N2016) );
  AO21X1 U651 ( .IN1(N50), .IN2(n481), .IN3(n593), .Q(n592) );
  XOR2X1 U652 ( .IN1(n594), .IN2(keyinput1), .Q(n593) );
  NAND2X0 U653 ( .IN1(N75), .IN2(n484), .QN(n594) );
  AO221X1 U654 ( .IN1(N63), .IN2(n480), .IN3(N51), .IN4(n481), .IN5(n595), .Q(
        N2014) );
  AO22X1 U655 ( .IN1(N89), .IN2(n483), .IN3(N76), .IN4(n484), .Q(n595) );
  AO221X1 U656 ( .IN1(N64), .IN2(n480), .IN3(N52), .IN4(n481), .IN5(n596), .Q(
        N2012) );
  AO22X1 U657 ( .IN1(N90), .IN2(n483), .IN3(N77), .IN4(n484), .Q(n596) );
  AO221X1 U658 ( .IN1(N65), .IN2(n480), .IN3(N53), .IN4(n481), .IN5(n597), .Q(
        N2010) );
  AO22X1 U659 ( .IN1(N91), .IN2(n483), .IN3(N78), .IN4(n484), .Q(n597) );
  AND2X1 U660 ( .IN1(N227), .IN2(N234), .Q(n484) );
  NOR2X0 U661 ( .IN1(N227), .IN2(N234), .QN(n483) );
  NOR2X0 U662 ( .IN1(n590), .IN2(N234), .QN(n481) );
  INVX0 U663 ( .INP(n589), .ZN(n480) );
  NAND2X0 U664 ( .IN1(N234), .IN2(n590), .QN(n589) );
  INVX0 U665 ( .INP(N227), .ZN(n590) );
  AOI22X1 U666 ( .IN1(N325), .IN2(n598), .IN3(N231), .IN4(n599), .QN(N1726) );
  INVX0 U667 ( .INP(N1277), .ZN(N1448) );
  NAND2X0 U668 ( .IN1(N325), .IN2(n600), .QN(N1269) );
  NOR2X0 U669 ( .IN1(n599), .IN2(n598), .QN(N1277) );
  NAND4X0 U670 ( .IN1(N44), .IN2(N132), .IN3(N82), .IN4(N96), .QN(n598) );
  NAND4X0 U671 ( .IN1(N69), .IN2(N120), .IN3(N57), .IN4(N108), .QN(n599) );
  NAND2X0 U672 ( .IN1(N231), .IN2(n600), .QN(N1029) );
  INVX0 U673 ( .INP(N1028), .ZN(n600) );
  NAND2X0 U674 ( .IN1(N7), .IN2(N237), .QN(N1028) );
  AND2X1 U675 ( .IN1(N94), .IN2(N219), .Q(N1026) );
endmodule

