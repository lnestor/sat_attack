
module c1355_NR1550 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, 
        G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, 
        G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
        G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, 
        G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, 
        G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, 
        G6, G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, 
        keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, 
        keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, 
        keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, 
        keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, 
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, 
        keyinput99, keyinput100, keyinput101, keyinput102, keyinput103, 
        keyinput104, keyinput105, keyinput106, keyinput107, keyinput108, 
        keyinput109, keyinput110, keyinput111, keyinput112, keyinput113, 
        keyinput114, keyinput115, keyinput116, keyinput117, keyinput118, 
        keyinput119, keyinput120, keyinput121, keyinput122, keyinput123, 
        keyinput124, keyinput125, keyinput126, keyinput127, keyinput128, 
        keyinput129, keyinput130, keyinput131, keyinput132, keyinput133, 
        keyinput134, keyinput135, keyinput136, keyinput137, keyinput138, 
        keyinput139, keyinput140, keyinput141, keyinput142, keyinput143, 
        keyinput144, keyinput145, keyinput146, keyinput147, keyinput148, 
        keyinput149, keyinput150, keyinput151, keyinput152, keyinput153, 
        keyinput154 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9,
         keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
         keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21,
         keyinput22, keyinput23, keyinput24, keyinput25,
         keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341;

  DELLN2X2 U657 ( .INP(keyinput16), .Z(n814) );
  DELLN2X2 U658 ( .INP(keyinput19), .Z(n815) );
  DELLN2X2 U659 ( .INP(keyinput20), .Z(n816) );
  DELLN2X2 U660 ( .INP(keyinput154), .Z(n817) );
  DELLN2X2 U661 ( .INP(keyinput152), .Z(n818) );
  DELLN2X2 U662 ( .INP(keyinput150), .Z(n819) );
  DELLN2X2 U663 ( .INP(keyinput149), .Z(n820) );
  DELLN2X2 U664 ( .INP(keyinput148), .Z(n821) );
  DELLN2X2 U665 ( .INP(keyinput147), .Z(n822) );
  DELLN2X2 U666 ( .INP(keyinput146), .Z(n823) );
  DELLN2X2 U667 ( .INP(keyinput145), .Z(n824) );
  DELLN2X2 U668 ( .INP(keyinput143), .Z(n825) );
  DELLN2X2 U669 ( .INP(keyinput142), .Z(n826) );
  DELLN2X2 U670 ( .INP(keyinput140), .Z(n827) );
  DELLN2X2 U671 ( .INP(keyinput139), .Z(n828) );
  DELLN2X2 U672 ( .INP(keyinput138), .Z(n829) );
  DELLN2X2 U673 ( .INP(keyinput137), .Z(n830) );
  DELLN2X2 U674 ( .INP(keyinput136), .Z(n831) );
  DELLN2X2 U675 ( .INP(keyinput134), .Z(n832) );
  DELLN2X2 U676 ( .INP(keyinput133), .Z(n833) );
  DELLN2X2 U677 ( .INP(keyinput132), .Z(n834) );
  DELLN2X2 U678 ( .INP(keyinput131), .Z(n835) );
  DELLN2X2 U679 ( .INP(keyinput130), .Z(n836) );
  DELLN2X2 U680 ( .INP(keyinput129), .Z(n837) );
  DELLN2X2 U681 ( .INP(keyinput128), .Z(n838) );
  DELLN2X2 U682 ( .INP(keyinput127), .Z(n839) );
  DELLN2X2 U683 ( .INP(keyinput126), .Z(n840) );
  DELLN2X2 U684 ( .INP(keyinput125), .Z(n841) );
  DELLN2X2 U685 ( .INP(keyinput124), .Z(n842) );
  DELLN2X2 U686 ( .INP(keyinput122), .Z(n843) );
  DELLN2X2 U687 ( .INP(keyinput121), .Z(n844) );
  DELLN2X2 U688 ( .INP(keyinput120), .Z(n845) );
  DELLN2X2 U689 ( .INP(keyinput119), .Z(n846) );
  DELLN2X2 U690 ( .INP(keyinput115), .Z(n847) );
  DELLN2X2 U691 ( .INP(keyinput114), .Z(n848) );
  DELLN2X2 U692 ( .INP(keyinput31), .Z(n849) );
  DELLN2X2 U693 ( .INP(keyinput30), .Z(n850) );
  DELLN2X2 U694 ( .INP(keyinput29), .Z(n851) );
  DELLN2X2 U695 ( .INP(keyinput28), .Z(n852) );
  DELLN2X2 U696 ( .INP(keyinput14), .Z(n853) );
  DELLN2X2 U697 ( .INP(keyinput7), .Z(n854) );
  DELLN2X2 U698 ( .INP(keyinput5), .Z(n855) );
  DELLN2X2 U699 ( .INP(keyinput151), .Z(n856) );
  DELLN2X2 U700 ( .INP(keyinput144), .Z(n857) );
  DELLN2X2 U701 ( .INP(keyinput141), .Z(n858) );
  DELLN2X2 U702 ( .INP(keyinput135), .Z(n859) );
  DELLN2X2 U703 ( .INP(keyinput123), .Z(n860) );
  DELLN2X2 U704 ( .INP(keyinput118), .Z(n861) );
  DELLN2X2 U705 ( .INP(keyinput117), .Z(n862) );
  DELLN2X2 U706 ( .INP(keyinput116), .Z(n863) );
  DELLN2X2 U707 ( .INP(keyinput153), .Z(n864) );
  DELLN2X2 U708 ( .INP(keyinput94), .Z(n865) );
  DELLN2X2 U709 ( .INP(keyinput91), .Z(n866) );
  DELLN2X2 U710 ( .INP(keyinput83), .Z(n867) );
  DELLN2X2 U711 ( .INP(keyinput82), .Z(n868) );
  DELLN2X2 U712 ( .INP(keyinput71), .Z(n869) );
  DELLN2X2 U713 ( .INP(keyinput69), .Z(n870) );
  DELLN2X2 U714 ( .INP(keyinput56), .Z(n871) );
  DELLN2X2 U715 ( .INP(keyinput53), .Z(n872) );
  DELLN2X2 U716 ( .INP(keyinput50), .Z(n873) );
  DELLN2X2 U717 ( .INP(keyinput47), .Z(n874) );
  DELLN2X2 U718 ( .INP(keyinput22), .Z(n875) );
  DELLN2X2 U719 ( .INP(keyinput104), .Z(n876) );
  DELLN2X2 U720 ( .INP(keyinput100), .Z(n877) );
  DELLN2X2 U721 ( .INP(keyinput93), .Z(n878) );
  DELLN2X2 U722 ( .INP(keyinput90), .Z(n879) );
  DELLN2X2 U723 ( .INP(keyinput87), .Z(n880) );
  DELLN2X2 U724 ( .INP(keyinput81), .Z(n881) );
  DELLN2X2 U725 ( .INP(keyinput57), .Z(n882) );
  DELLN2X2 U726 ( .INP(keyinput55), .Z(n883) );
  DELLN2X2 U727 ( .INP(keyinput43), .Z(n884) );
  DELLN2X2 U728 ( .INP(keyinput36), .Z(n885) );
  DELLN2X2 U729 ( .INP(keyinput33), .Z(n886) );
  DELLN2X2 U730 ( .INP(keyinput27), .Z(n887) );
  DELLN2X2 U731 ( .INP(keyinput26), .Z(n888) );
  DELLN2X2 U732 ( .INP(keyinput21), .Z(n889) );
  DELLN2X2 U733 ( .INP(keyinput15), .Z(n890) );
  DELLN2X2 U734 ( .INP(keyinput13), .Z(n891) );
  DELLN2X2 U735 ( .INP(keyinput11), .Z(n892) );
  DELLN2X2 U736 ( .INP(keyinput9), .Z(n893) );
  DELLN2X2 U737 ( .INP(keyinput4), .Z(n894) );
  DELLN2X2 U738 ( .INP(keyinput0), .Z(n895) );
  DELLN2X2 U739 ( .INP(keyinput113), .Z(n896) );
  DELLN2X2 U740 ( .INP(keyinput111), .Z(n897) );
  DELLN2X2 U741 ( .INP(keyinput110), .Z(n898) );
  DELLN2X2 U742 ( .INP(keyinput109), .Z(n899) );
  DELLN2X2 U743 ( .INP(keyinput108), .Z(n900) );
  DELLN2X2 U744 ( .INP(keyinput107), .Z(n901) );
  DELLN2X2 U745 ( .INP(keyinput105), .Z(n902) );
  DELLN2X2 U746 ( .INP(keyinput99), .Z(n903) );
  DELLN2X2 U747 ( .INP(keyinput98), .Z(n904) );
  DELLN2X2 U748 ( .INP(keyinput96), .Z(n905) );
  DELLN2X2 U749 ( .INP(keyinput95), .Z(n906) );
  DELLN2X2 U750 ( .INP(keyinput92), .Z(n907) );
  DELLN2X2 U751 ( .INP(keyinput88), .Z(n908) );
  DELLN2X2 U752 ( .INP(keyinput84), .Z(n909) );
  DELLN2X2 U753 ( .INP(keyinput78), .Z(n910) );
  DELLN2X2 U754 ( .INP(keyinput76), .Z(n911) );
  DELLN2X2 U755 ( .INP(keyinput75), .Z(n912) );
  DELLN2X2 U756 ( .INP(keyinput73), .Z(n913) );
  DELLN2X2 U757 ( .INP(keyinput72), .Z(n914) );
  DELLN2X2 U758 ( .INP(keyinput70), .Z(n915) );
  DELLN2X2 U759 ( .INP(keyinput68), .Z(n916) );
  DELLN2X2 U760 ( .INP(keyinput67), .Z(n917) );
  DELLN2X2 U761 ( .INP(keyinput66), .Z(n918) );
  DELLN2X2 U762 ( .INP(keyinput63), .Z(n919) );
  DELLN2X2 U763 ( .INP(keyinput61), .Z(n920) );
  DELLN2X2 U764 ( .INP(keyinput54), .Z(n921) );
  DELLN2X2 U765 ( .INP(keyinput51), .Z(n922) );
  DELLN2X2 U766 ( .INP(keyinput49), .Z(n923) );
  DELLN2X2 U767 ( .INP(keyinput46), .Z(n924) );
  DELLN2X2 U768 ( .INP(keyinput35), .Z(n925) );
  DELLN2X2 U769 ( .INP(keyinput32), .Z(n926) );
  DELLN2X2 U770 ( .INP(keyinput6), .Z(n927) );
  DELLN2X2 U771 ( .INP(keyinput112), .Z(n928) );
  DELLN2X2 U772 ( .INP(keyinput101), .Z(n929) );
  DELLN2X2 U773 ( .INP(keyinput97), .Z(n930) );
  DELLN2X2 U774 ( .INP(keyinput79), .Z(n931) );
  DELLN2X2 U775 ( .INP(keyinput60), .Z(n932) );
  DELLN2X2 U776 ( .INP(keyinput45), .Z(n933) );
  DELLN2X2 U777 ( .INP(keyinput41), .Z(n934) );
  DELLN2X2 U778 ( .INP(keyinput38), .Z(n935) );
  DELLN2X2 U779 ( .INP(keyinput106), .Z(n936) );
  DELLN2X2 U780 ( .INP(keyinput103), .Z(n937) );
  DELLN2X2 U781 ( .INP(keyinput102), .Z(n938) );
  DELLN2X2 U782 ( .INP(keyinput89), .Z(n939) );
  DELLN2X2 U783 ( .INP(keyinput86), .Z(n940) );
  DELLN2X2 U784 ( .INP(keyinput85), .Z(n941) );
  DELLN2X2 U785 ( .INP(keyinput80), .Z(n942) );
  DELLN2X2 U786 ( .INP(keyinput77), .Z(n943) );
  DELLN2X2 U787 ( .INP(keyinput74), .Z(n944) );
  DELLN2X2 U788 ( .INP(keyinput65), .Z(n945) );
  DELLN2X2 U789 ( .INP(keyinput64), .Z(n946) );
  DELLN2X2 U790 ( .INP(keyinput62), .Z(n947) );
  DELLN2X2 U791 ( .INP(keyinput59), .Z(n948) );
  DELLN2X2 U792 ( .INP(keyinput58), .Z(n949) );
  DELLN2X2 U793 ( .INP(keyinput52), .Z(n950) );
  DELLN2X2 U794 ( .INP(keyinput48), .Z(n951) );
  DELLN2X2 U795 ( .INP(keyinput44), .Z(n952) );
  DELLN2X2 U796 ( .INP(keyinput42), .Z(n953) );
  DELLN2X2 U797 ( .INP(keyinput40), .Z(n954) );
  DELLN2X2 U798 ( .INP(keyinput39), .Z(n955) );
  DELLN2X2 U799 ( .INP(keyinput37), .Z(n956) );
  DELLN2X2 U800 ( .INP(keyinput34), .Z(n957) );
  DELLN2X2 U801 ( .INP(keyinput25), .Z(n958) );
  DELLN2X2 U802 ( .INP(keyinput24), .Z(n959) );
  DELLN2X2 U803 ( .INP(keyinput18), .Z(n960) );
  DELLN2X2 U804 ( .INP(keyinput12), .Z(n961) );
  DELLN2X2 U805 ( .INP(keyinput10), .Z(n962) );
  DELLN2X2 U806 ( .INP(keyinput8), .Z(n963) );
  DELLN2X2 U807 ( .INP(keyinput3), .Z(n964) );
  DELLN2X2 U808 ( .INP(keyinput2), .Z(n965) );
  DELLN2X2 U809 ( .INP(keyinput1), .Z(n966) );
  INVX0 U810 ( .INP(n968), .ZN(n967) );
  DELLN2X2 U811 ( .INP(keyinput23), .Z(n968) );
  DELLN2X2 U812 ( .INP(keyinput17), .Z(n969) );
  DELLN2X2 U813 ( .INP(G37), .Z(n970) );
  DELLN2X2 U814 ( .INP(G14), .Z(n971) );
  DELLN2X2 U815 ( .INP(G20), .Z(n972) );
  DELLN2X2 U816 ( .INP(G34), .Z(n973) );
  INVX0 U817 ( .INP(n975), .ZN(n974) );
  DELLN2X2 U818 ( .INP(G33), .Z(n975) );
  INVX0 U819 ( .INP(n977), .ZN(n976) );
  DELLN2X2 U820 ( .INP(G38), .Z(n977) );
  DELLN2X2 U821 ( .INP(G31), .Z(n978) );
  DELLN2X2 U822 ( .INP(G30), .Z(n979) );
  DELLN2X2 U823 ( .INP(G13), .Z(n980) );
  DELLN2X2 U824 ( .INP(G9), .Z(n981) );
  DELLN2X2 U825 ( .INP(G39), .Z(n982) );
  DELLN2X2 U826 ( .INP(G36), .Z(n983) );
  DELLN2X2 U827 ( .INP(G35), .Z(n984) );
  DELLN2X2 U828 ( .INP(G40), .Z(n985) );
  INVX0 U829 ( .INP(n987), .ZN(n986) );
  DELLN2X2 U830 ( .INP(G19), .Z(n987) );
  DELLN2X2 U831 ( .INP(G1), .Z(n988) );
  DELLN2X2 U832 ( .INP(G10), .Z(n989) );
  INVX0 U833 ( .INP(n991), .ZN(n990) );
  DELLN2X2 U834 ( .INP(G23), .Z(n991) );
  INVX0 U835 ( .INP(n993), .ZN(n992) );
  DELLN2X2 U836 ( .INP(G26), .Z(n993) );
  DELLN2X2 U837 ( .INP(G2), .Z(n994) );
  INVX0 U838 ( .INP(n996), .ZN(n995) );
  DELLN2X2 U839 ( .INP(G3), .Z(n996) );
  INVX0 U840 ( .INP(n998), .ZN(n997) );
  DELLN2X2 U841 ( .INP(G28), .Z(n998) );
  INVX0 U842 ( .INP(n1000), .ZN(n999) );
  DELLN2X2 U843 ( .INP(G16), .Z(n1000) );
  INVX0 U844 ( .INP(n1002), .ZN(n1001) );
  DELLN2X2 U845 ( .INP(G4), .Z(n1002) );
  DELLN2X2 U846 ( .INP(G21), .Z(n1003) );
  DELLN2X2 U847 ( .INP(G11), .Z(n1004) );
  INVX0 U848 ( .INP(n1006), .ZN(n1005) );
  DELLN2X2 U849 ( .INP(G32), .Z(n1006) );
  INVX0 U850 ( .INP(n1008), .ZN(n1007) );
  DELLN2X2 U851 ( .INP(G5), .Z(n1008) );
  DELLN2X2 U852 ( .INP(G15), .Z(n1009) );
  INVX0 U853 ( .INP(n1011), .ZN(n1010) );
  DELLN2X2 U854 ( .INP(G17), .Z(n1011) );
  DELLN2X2 U855 ( .INP(G12), .Z(n1012) );
  DELLN2X2 U856 ( .INP(G18), .Z(n1013) );
  DELLN2X2 U857 ( .INP(G7), .Z(n1014) );
  DELLN2X2 U858 ( .INP(G24), .Z(n1015) );
  DELLN2X2 U859 ( .INP(G22), .Z(n1016) );
  DELLN2X2 U860 ( .INP(G27), .Z(n1017) );
  DELLN2X2 U861 ( .INP(G8), .Z(n1018) );
  DELLN2X2 U862 ( .INP(G6), .Z(n1019) );
  DELLN2X2 U863 ( .INP(G29), .Z(n1020) );
  INVX0 U864 ( .INP(n1022), .ZN(n1021) );
  DELLN2X2 U865 ( .INP(G41), .Z(n1022) );
  DELLN2X2 U866 ( .INP(G25), .Z(n1023) );
  AO21X1 U867 ( .IN1(n1005), .IN2(n967), .IN3(n1024), .Q(G1355) );
  XOR2X1 U868 ( .IN1(n1025), .IN2(n1026), .Q(n1024) );
  NOR2X0 U869 ( .IN1(n1027), .IN2(n1028), .QN(n1026) );
  NAND2X0 U870 ( .IN1(n968), .IN2(n1006), .QN(n1025) );
  XOR2X1 U871 ( .IN1(n1029), .IN2(n1030), .Q(G1353) );
  NOR2X0 U872 ( .IN1(n1031), .IN2(n1028), .QN(n1030) );
  NOR2X0 U873 ( .IN1(n1032), .IN2(n1033), .QN(G1352) );
  XOR2X1 U874 ( .IN1(n1034), .IN2(n887), .Q(n1033) );
  OR3X1 U875 ( .IN1(n1035), .IN2(n1020), .IN3(n1028), .Q(n1034) );
  OA21X1 U876 ( .IN1(n1035), .IN2(n1028), .IN3(n1020), .Q(n1032) );
  XOR2X1 U877 ( .IN1(n1036), .IN2(n998), .Q(G1351) );
  NAND2X0 U878 ( .IN1(n1037), .IN2(n1038), .QN(n1036) );
  XOR2X1 U879 ( .IN1(n1039), .IN2(n1017), .Q(G1350) );
  NAND2X0 U880 ( .IN1(n1037), .IN2(n1040), .QN(n1039) );
  XOR2X1 U881 ( .IN1(n1041), .IN2(n993), .Q(G1349) );
  NAND2X0 U882 ( .IN1(n1037), .IN2(n1042), .QN(n1041) );
  XOR2X1 U883 ( .IN1(n1043), .IN2(n1023), .Q(G1348) );
  NAND2X0 U884 ( .IN1(n1037), .IN2(n1044), .QN(n1043) );
  AND3X1 U885 ( .IN1(n1045), .IN2(n1046), .IN3(n1047), .Q(n1037) );
  OA21X1 U886 ( .IN1(n1048), .IN2(n990), .IN3(n1049), .Q(G1346) );
  XOR2X1 U887 ( .IN1(n1050), .IN2(n888), .Q(n1049) );
  NAND3X0 U888 ( .IN1(n1040), .IN2(n990), .IN3(n1051), .QN(n1050) );
  NOR2X0 U889 ( .IN1(n1052), .IN2(n1053), .QN(n1048) );
  XOR2X1 U890 ( .IN1(n1054), .IN2(n1016), .Q(G1345) );
  NAND2X0 U891 ( .IN1(n1051), .IN2(n1042), .QN(n1054) );
  XOR2X1 U892 ( .IN1(n1055), .IN2(n1003), .Q(G1344) );
  NAND2X0 U893 ( .IN1(n1051), .IN2(n1044), .QN(n1055) );
  INVX0 U894 ( .INP(n1053), .ZN(n1051) );
  XOR2X1 U895 ( .IN1(n1056), .IN2(n1057), .Q(G1343) );
  NOR2X0 U896 ( .IN1(n1027), .IN2(n1058), .QN(n1057) );
  XOR2X1 U897 ( .IN1(n986), .IN2(n1059), .Q(G1342) );
  NOR2X0 U898 ( .IN1(n1052), .IN2(n1058), .QN(n1059) );
  XNOR2X1 U899 ( .IN1(n1013), .IN2(n1060), .Q(G1341) );
  NOR2X0 U900 ( .IN1(n1031), .IN2(n1058), .QN(n1060) );
  XOR2X1 U901 ( .IN1(n1010), .IN2(n1061), .Q(G1340) );
  NOR2X0 U902 ( .IN1(n1035), .IN2(n1058), .QN(n1061) );
  NAND3X0 U903 ( .IN1(n1047), .IN2(n1062), .IN3(n1063), .QN(n1058) );
  AND3X1 U904 ( .IN1(n1064), .IN2(n1065), .IN3(n1066), .Q(n1047) );
  XOR2X1 U905 ( .IN1(n999), .IN2(n1067), .Q(G1339) );
  NOR2X0 U906 ( .IN1(n1064), .IN2(n1068), .QN(n1067) );
  XNOR2X1 U907 ( .IN1(n1009), .IN2(n1069), .Q(G1338) );
  NOR2X0 U908 ( .IN1(n1070), .IN2(n1068), .QN(n1069) );
  XOR2X1 U909 ( .IN1(n1071), .IN2(n1072), .Q(G1337) );
  NOR2X0 U910 ( .IN1(n1062), .IN2(n1068), .QN(n1072) );
  XOR2X1 U911 ( .IN1(n1073), .IN2(n1074), .Q(G1336) );
  NOR2X0 U912 ( .IN1(n1046), .IN2(n1068), .QN(n1074) );
  NAND3X0 U913 ( .IN1(n1035), .IN2(n1042), .IN3(n1075), .QN(n1068) );
  XNOR2X1 U914 ( .IN1(n1012), .IN2(n1076), .Q(G1335) );
  NOR2X0 U915 ( .IN1(n1064), .IN2(n1077), .QN(n1076) );
  XNOR2X1 U916 ( .IN1(n1004), .IN2(n1078), .Q(G1334) );
  NOR2X0 U917 ( .IN1(n1070), .IN2(n1077), .QN(n1078) );
  XOR2X1 U918 ( .IN1(n1079), .IN2(n1080), .Q(G1333) );
  NOR2X0 U919 ( .IN1(n1062), .IN2(n1077), .QN(n1080) );
  XOR2X1 U920 ( .IN1(n1081), .IN2(n1018), .Q(G1331) );
  NAND2X0 U921 ( .IN1(n1082), .IN2(n1083), .QN(n1081) );
  XOR2X1 U922 ( .IN1(n1084), .IN2(n1014), .Q(G1330) );
  NAND2X0 U923 ( .IN1(n1082), .IN2(n1066), .QN(n1084) );
  XOR2X1 U924 ( .IN1(n1085), .IN2(n1008), .Q(G1328) );
  NAND2X0 U925 ( .IN1(n1082), .IN2(n1063), .QN(n1085) );
  XOR2X1 U926 ( .IN1(n1001), .IN2(n1086), .Q(G1327) );
  NOR2X0 U927 ( .IN1(n1064), .IN2(n1087), .QN(n1086) );
  NOR2X0 U928 ( .IN1(n1088), .IN2(n1089), .QN(G1326) );
  XOR2X1 U929 ( .IN1(n958), .IN2(n1090), .Q(n1089) );
  NOR2X0 U930 ( .IN1(n1091), .IN2(n995), .QN(n1090) );
  NOR3X0 U931 ( .IN1(n1087), .IN2(n1091), .IN3(n1070), .QN(n1088) );
  NOR3X0 U932 ( .IN1(n1070), .IN2(n995), .IN3(n1087), .QN(n1091) );
  OA21X1 U933 ( .IN1(n1092), .IN2(n1093), .IN3(n1094), .Q(G1325) );
  XOR2X1 U934 ( .IN1(n959), .IN2(n1095), .Q(n1094) );
  NOR2X0 U935 ( .IN1(n1096), .IN2(n1093), .QN(n1095) );
  XNOR2X1 U936 ( .IN1(n1097), .IN2(n875), .Q(n1093) );
  OR2X1 U937 ( .IN1(n1096), .IN2(n1092), .Q(n1097) );
  NAND2X0 U938 ( .IN1(n1098), .IN2(n1045), .QN(n1096) );
  XOR3X1 U939 ( .IN1(n849), .IN2(n978), .IN3(n1099), .Q(G1354) );
  NOR2X0 U940 ( .IN1(n1052), .IN2(n1028), .QN(n1099) );
  NAND4X0 U941 ( .IN1(n1046), .IN2(n1065), .IN3(n1070), .IN4(n1100), .QN(n1028) );
  NOR2X0 U942 ( .IN1(n1064), .IN2(n1062), .QN(n1100) );
  XOR3X1 U943 ( .IN1(n850), .IN2(n981), .IN3(n1101), .Q(G1332) );
  NOR2X0 U944 ( .IN1(n1046), .IN2(n1077), .QN(n1101) );
  NAND3X0 U945 ( .IN1(n1035), .IN2(n1042), .IN3(n1102), .QN(n1077) );
  XOR3X1 U946 ( .IN1(n817), .IN2(n1015), .IN3(n1103), .Q(G1347) );
  XOR2X1 U947 ( .IN1(n1104), .IN2(n1105), .Q(n1103) );
  NOR2X0 U948 ( .IN1(n1027), .IN2(n1053), .QN(n1105) );
  NAND4X0 U949 ( .IN1(n1106), .IN2(n1062), .IN3(n1070), .IN4(n1065), .QN(n1053) );
  NAND2X0 U950 ( .IN1(n1107), .IN2(n1108), .QN(n1065) );
  NAND3X0 U951 ( .IN1(n1027), .IN2(n1109), .IN3(n1052), .QN(n1108) );
  XOR2X1 U952 ( .IN1(n1110), .IN2(n1042), .Q(n1109) );
  INVX0 U953 ( .INP(n1031), .ZN(n1042) );
  NOR2X0 U954 ( .IN1(n1035), .IN2(n816), .QN(n1110) );
  NAND3X0 U955 ( .IN1(n1031), .IN2(n1111), .IN3(n1035), .QN(n1107) );
  INVX0 U956 ( .INP(n1044), .ZN(n1035) );
  XOR2X1 U957 ( .IN1(n1112), .IN2(n1038), .Q(n1111) );
  NOR2X0 U958 ( .IN1(n815), .IN2(n1052), .QN(n1112) );
  NAND2X0 U959 ( .IN1(n1113), .IN2(n1114), .QN(n1104) );
  NAND4X0 U960 ( .IN1(n1115), .IN2(n1116), .IN3(n1117), .IN4(n1118), .QN(n1114) );
  NOR4X0 U961 ( .IN1(n1119), .IN2(n1120), .IN3(n1121), .IN4(n1122), .QN(n1118)
         );
  XOR3X1 U962 ( .IN1(n823), .IN2(n901), .IN3(n1073), .Q(n1122) );
  XOR3X1 U963 ( .IN1(n824), .IN2(n902), .IN3(n1021), .Q(n1121) );
  NAND3X0 U964 ( .IN1(n1123), .IN2(n1124), .IN3(n1125), .QN(n1120) );
  XOR3X1 U965 ( .IN1(n827), .IN2(n905), .IN3(n993), .Q(n1125) );
  XOR3X1 U966 ( .IN1(n826), .IN2(n904), .IN3(n971), .Q(n1124) );
  XOR3X1 U967 ( .IN1(n828), .IN2(n906), .IN3(n1023), .Q(n1123) );
  NAND4X0 U968 ( .IN1(n1126), .IN2(n1127), .IN3(n1128), .IN4(n1129), .QN(n1119) );
  NOR3X0 U969 ( .IN1(n1130), .IN2(n1131), .IN3(n1132), .QN(n1129) );
  XOR3X1 U970 ( .IN1(n833), .IN2(n911), .IN3(n1133), .Q(n1132) );
  XNOR3X1 U971 ( .IN1(n859), .IN2(n931), .IN3(n982), .Q(n1131) );
  XOR3X1 U972 ( .IN1(n832), .IN2(n910), .IN3(n1134), .Q(n1130) );
  XOR3X1 U973 ( .IN1(n830), .IN2(n908), .IN3(n973), .Q(n1128) );
  XOR3X1 U974 ( .IN1(n829), .IN2(n907), .IN3(n987), .Q(n1127) );
  XOR3X1 U975 ( .IN1(n831), .IN2(n909), .IN3(n991), .Q(n1126) );
  NOR4X0 U976 ( .IN1(n1135), .IN2(n1136), .IN3(n1137), .IN4(n1138), .QN(n1117)
         );
  XOR3X1 U977 ( .IN1(n818), .IN2(n896), .IN3(n1029), .Q(n1138) );
  XNOR3X1 U978 ( .IN1(n856), .IN2(n928), .IN3(n1009), .Q(n1137) );
  NAND3X0 U979 ( .IN1(n1139), .IN2(n1140), .IN3(n1141), .QN(n1136) );
  XOR3X1 U980 ( .IN1(n820), .IN2(n898), .IN3(n1015), .Q(n1141) );
  XOR3X1 U981 ( .IN1(n819), .IN2(n897), .IN3(n1018), .Q(n1140) );
  XOR3X1 U982 ( .IN1(n822), .IN2(n900), .IN3(n996), .Q(n1139) );
  NAND4X0 U983 ( .IN1(n1142), .IN2(n1143), .IN3(n1144), .IN4(n1145), .QN(n1135) );
  NOR2X0 U984 ( .IN1(n1146), .IN2(n1147), .QN(n1145) );
  XOR2X1 U985 ( .IN1(n974), .IN2(n879), .Q(n1147) );
  XOR2X1 U986 ( .IN1(n997), .IN2(n876), .Q(n1146) );
  XOR2X1 U987 ( .IN1(n941), .IN2(n1011), .Q(n1144) );
  XOR2X1 U988 ( .IN1(n938), .IN2(n972), .Q(n1143) );
  XOR2X1 U989 ( .IN1(n939), .IN2(n1000), .Q(n1142) );
  NOR4X0 U990 ( .IN1(n1148), .IN2(n1149), .IN3(n1150), .IN4(n1151), .QN(n1116)
         );
  XOR2X1 U991 ( .IN1(n940), .IN2(n1012), .Q(n1151) );
  XOR3X1 U992 ( .IN1(n821), .IN2(n899), .IN3(n1013), .Q(n1150) );
  NAND3X0 U993 ( .IN1(n1152), .IN2(n1153), .IN3(n1154), .QN(n1149) );
  XOR3X1 U994 ( .IN1(n825), .IN2(n903), .IN3(n1079), .Q(n1154) );
  XNOR3X1 U995 ( .IN1(n857), .IN2(n929), .IN3(n970), .Q(n1153) );
  XNOR3X1 U996 ( .IN1(n858), .IN2(n930), .IN3(n1004), .Q(n1152) );
  NAND4X0 U997 ( .IN1(n1155), .IN2(n1156), .IN3(n1157), .IN4(n1158), .QN(n1148) );
  XOR2X1 U998 ( .IN1(n944), .IN2(n977), .Q(n1158) );
  NOR2X0 U999 ( .IN1(n1159), .IN2(n1160), .QN(n1157) );
  XNOR2X1 U1000 ( .IN1(n983), .IN2(n866), .Q(n1160) );
  XNOR2X1 U1001 ( .IN1(n985), .IN2(n868), .Q(n1159) );
  XOR3X1 U1002 ( .IN1(n835), .IN2(n913), .IN3(n1161), .Q(n1156) );
  XOR3X1 U1003 ( .IN1(n834), .IN2(n912), .IN3(n1162), .Q(n1155) );
  NOR4X0 U1004 ( .IN1(n1163), .IN2(n1164), .IN3(n1165), .IN4(n1166), .QN(n1115) );
  XOR2X1 U1005 ( .IN1(n942), .IN2(n1014), .Q(n1166) );
  XOR2X1 U1006 ( .IN1(n936), .IN2(n1019), .Q(n1165) );
  NAND3X0 U1007 ( .IN1(n1167), .IN2(n1168), .IN3(n1169), .QN(n1164) );
  XOR2X1 U1008 ( .IN1(n1001), .IN2(n877), .Q(n1169) );
  XOR2X1 U1009 ( .IN1(n1007), .IN2(n881), .Q(n1168) );
  XNOR2X1 U1010 ( .IN1(n984), .IN2(n865), .Q(n1167) );
  NAND4X0 U1011 ( .IN1(n1170), .IN2(n1171), .IN3(n1172), .IN4(n1173), .QN(
        n1163) );
  XNOR2X1 U1012 ( .IN1(n1016), .IN2(n867), .Q(n1173) );
  NOR2X0 U1013 ( .IN1(n1174), .IN2(n1175), .QN(n1172) );
  XOR2X1 U1014 ( .IN1(n943), .IN2(n994), .Q(n1175) );
  XOR2X1 U1015 ( .IN1(n937), .IN2(n1017), .Q(n1174) );
  XOR2X1 U1016 ( .IN1(n1176), .IN2(n880), .Q(n1171) );
  XOR2X1 U1017 ( .IN1(n1005), .IN2(n878), .Q(n1170) );
  XNOR2X1 U1018 ( .IN1(n1177), .IN2(n864), .Q(n1113) );
  NAND4X0 U1019 ( .IN1(n1178), .IN2(n1179), .IN3(n1180), .IN4(n1181), .QN(
        n1177) );
  NOR4X0 U1020 ( .IN1(n1182), .IN2(n1183), .IN3(n1184), .IN4(n1185), .QN(n1181) );
  XNOR3X1 U1021 ( .IN1(n862), .IN2(n934), .IN3(n985), .Q(n1185) );
  XNOR3X1 U1022 ( .IN1(n863), .IN2(n935), .IN3(n982), .Q(n1184) );
  NAND3X0 U1023 ( .IN1(n1186), .IN2(n1187), .IN3(n1188), .QN(n1183) );
  XOR3X1 U1024 ( .IN1(n837), .IN2(n915), .IN3(n1018), .Q(n1188) );
  XOR3X1 U1025 ( .IN1(n836), .IN2(n914), .IN3(n979), .Q(n1187) );
  XOR3X1 U1026 ( .IN1(n838), .IN2(n916), .IN3(n1013), .Q(n1186) );
  NAND4X0 U1027 ( .IN1(n1189), .IN2(n1190), .IN3(n1191), .IN4(n1192), .QN(
        n1182) );
  NOR3X0 U1028 ( .IN1(n1193), .IN2(n1194), .IN3(n1195), .QN(n1192) );
  XOR3X1 U1029 ( .IN1(n848), .IN2(n926), .IN3(n1161), .Q(n1195) );
  XOR3X1 U1030 ( .IN1(n842), .IN2(n920), .IN3(n1056), .Q(n1194) );
  XOR3X1 U1031 ( .IN1(n847), .IN2(n925), .IN3(n1133), .Q(n1193) );
  XOR3X1 U1032 ( .IN1(n840), .IN2(n918), .IN3(n980), .Q(n1191) );
  XOR3X1 U1033 ( .IN1(n839), .IN2(n917), .IN3(n996), .Q(n1190) );
  XOR3X1 U1034 ( .IN1(n841), .IN2(n919), .IN3(n998), .Q(n1189) );
  NOR4X0 U1035 ( .IN1(n1196), .IN2(n1197), .IN3(n1198), .IN4(n1199), .QN(n1180) );
  XNOR2X1 U1036 ( .IN1(n1015), .IN2(n870), .Q(n1199) );
  XOR2X1 U1037 ( .IN1(n990), .IN2(n884), .Q(n1198) );
  NAND3X0 U1038 ( .IN1(n1200), .IN2(n1201), .IN3(n1202), .QN(n1197) );
  XOR2X1 U1039 ( .IN1(n952), .IN2(n1011), .Q(n1202) );
  XOR2X1 U1040 ( .IN1(n953), .IN2(n1016), .Q(n1201) );
  XOR2X1 U1041 ( .IN1(n951), .IN2(n1000), .Q(n1200) );
  NAND4X0 U1042 ( .IN1(n1203), .IN2(n1204), .IN3(n1205), .IN4(n1206), .QN(
        n1196) );
  NOR2X0 U1043 ( .IN1(n1207), .IN2(n1208), .QN(n1206) );
  XNOR2X1 U1044 ( .IN1(n1009), .IN2(n869), .Q(n1208) );
  XNOR2X1 U1045 ( .IN1(n1004), .IN2(n871), .Q(n1207) );
  XOR2X1 U1046 ( .IN1(n956), .IN2(n988), .Q(n1205) );
  XOR2X1 U1047 ( .IN1(n949), .IN2(n989), .Q(n1204) );
  XOR3X1 U1048 ( .IN1(n843), .IN2(n921), .IN3(n1023), .Q(n1203) );
  NOR4X0 U1049 ( .IN1(n1209), .IN2(n1210), .IN3(n1211), .IN4(n1212), .QN(n1179) );
  XOR3X1 U1050 ( .IN1(n844), .IN2(n922), .IN3(n987), .Q(n1212) );
  XOR3X1 U1051 ( .IN1(n845), .IN2(n923), .IN3(n975), .Q(n1211) );
  NAND3X0 U1052 ( .IN1(n1213), .IN2(n1214), .IN3(n1215), .QN(n1210) );
  XNOR3X1 U1053 ( .IN1(n861), .IN2(n933), .IN3(n1012), .Q(n1215) );
  XOR2X1 U1054 ( .IN1(n955), .IN2(n1014), .Q(n1214) );
  XOR3X1 U1055 ( .IN1(n846), .IN2(n924), .IN3(n1176), .Q(n1213) );
  NAND4X0 U1056 ( .IN1(n1216), .IN2(n1217), .IN3(n1218), .IN4(n1219), .QN(
        n1209) );
  XOR2X1 U1057 ( .IN1(n950), .IN2(n1006), .Q(n1219) );
  NOR2X0 U1058 ( .IN1(n1220), .IN2(n1221), .QN(n1218) );
  XOR2X1 U1059 ( .IN1(n992), .IN2(n883), .Q(n1221) );
  XNOR2X1 U1060 ( .IN1(n983), .IN2(n873), .Q(n1220) );
  XOR2X1 U1061 ( .IN1(n948), .IN2(n1002), .Q(n1217) );
  XOR2X1 U1062 ( .IN1(n954), .IN2(n1008), .Q(n1216) );
  NOR4X0 U1063 ( .IN1(n1222), .IN2(n1223), .IN3(n1224), .IN4(n1225), .QN(n1178) );
  XOR2X1 U1064 ( .IN1(n945), .IN2(n1019), .Q(n1225) );
  XOR2X1 U1065 ( .IN1(n946), .IN2(n1022), .Q(n1224) );
  NAND3X0 U1066 ( .IN1(n1226), .IN2(n1227), .IN3(n1228), .QN(n1223) );
  XNOR2X1 U1067 ( .IN1(n984), .IN2(n872), .Q(n1228) );
  XOR2X1 U1068 ( .IN1(n976), .IN2(n886), .Q(n1227) );
  XNOR2X1 U1069 ( .IN1(n973), .IN2(n874), .Q(n1226) );
  NAND4X0 U1070 ( .IN1(n1229), .IN2(n1230), .IN3(n1231), .IN4(n1232), .QN(
        n1222) );
  NOR2X0 U1071 ( .IN1(n1233), .IN2(n1234), .QN(n1232) );
  XOR2X1 U1072 ( .IN1(n957), .IN2(n1020), .Q(n1234) );
  XOR2X1 U1073 ( .IN1(n947), .IN2(n1017), .Q(n1233) );
  XOR2X1 U1074 ( .IN1(n1071), .IN2(n882), .Q(n1231) );
  XOR2X1 U1075 ( .IN1(n1092), .IN2(n885), .Q(n1230) );
  XNOR3X1 U1076 ( .IN1(n860), .IN2(n932), .IN3(n970), .Q(n1229) );
  XOR3X1 U1077 ( .IN1(n851), .IN2(n1019), .IN3(n1235), .Q(G1329) );
  NAND2X0 U1078 ( .IN1(n1082), .IN2(n1045), .QN(n1235) );
  XOR2X1 U1079 ( .IN1(n1236), .IN2(n889), .Q(n1082) );
  NAND3X0 U1080 ( .IN1(n1031), .IN2(n1044), .IN3(n1075), .QN(n1236) );
  AND3X1 U1081 ( .IN1(n1038), .IN2(n1237), .IN3(n1052), .Q(n1075) );
  INVX0 U1082 ( .INP(n1027), .ZN(n1038) );
  XOR3X1 U1083 ( .IN1(n852), .IN2(n988), .IN3(n1238), .Q(G1324) );
  NAND2X0 U1084 ( .IN1(n1098), .IN2(n1063), .QN(n1238) );
  INVX0 U1085 ( .INP(n1087), .ZN(n1098) );
  NAND3X0 U1086 ( .IN1(n1031), .IN2(n1044), .IN3(n1102), .QN(n1087) );
  AND3X1 U1087 ( .IN1(n1040), .IN2(n1237), .IN3(n1027), .Q(n1102) );
  XOR3X1 U1088 ( .IN1(n1239), .IN2(n1240), .IN3(n1056), .Q(n1027) );
  XOR3X1 U1089 ( .IN1(n1006), .IN2(n998), .IN3(n1015), .Q(n1240) );
  OA21X1 U1090 ( .IN1(n1241), .IN2(n1242), .IN3(n1243), .Q(n1239) );
  NAND3X0 U1091 ( .IN1(n1022), .IN2(n1242), .IN3(n985), .QN(n1243) );
  XOR2X1 U1092 ( .IN1(n1244), .IN2(n1245), .Q(n1242) );
  INVX0 U1093 ( .INP(n1246), .ZN(n1244) );
  AND2X1 U1094 ( .IN1(n1022), .IN2(n985), .Q(n1241) );
  OAI21X1 U1095 ( .IN1(n1247), .IN2(n1045), .IN3(n1248), .QN(n1237) );
  NAND3X0 U1096 ( .IN1(n1249), .IN2(n1070), .IN3(n1250), .QN(n1248) );
  MUX21X1 U1097 ( .IN1(n1251), .IN2(n969), .S(n1046), .Q(n1250) );
  NOR2X0 U1098 ( .IN1(n969), .IN2(n1062), .QN(n1251) );
  INVX0 U1099 ( .INP(n1045), .ZN(n1062) );
  INVX0 U1100 ( .INP(n1066), .ZN(n1070) );
  XOR2X1 U1101 ( .IN1(n960), .IN2(n1083), .Q(n1249) );
  XNOR3X1 U1102 ( .IN1(n1252), .IN2(n1253), .IN3(n1254), .Q(n1045) );
  XOR2X1 U1103 ( .IN1(n1255), .IN2(n1256), .Q(n1254) );
  OA21X1 U1104 ( .IN1(n1257), .IN2(n1258), .IN3(n1259), .Q(n1256) );
  XOR2X1 U1105 ( .IN1(n961), .IN2(n1260), .Q(n1259) );
  NOR2X0 U1106 ( .IN1(n1257), .IN2(n1261), .QN(n1260) );
  INVX0 U1107 ( .INP(n1262), .ZN(n1261) );
  XOR2X1 U1108 ( .IN1(n1092), .IN2(n1019), .Q(n1258) );
  INVX0 U1109 ( .INP(n994), .ZN(n1092) );
  AND2X1 U1110 ( .IN1(n1263), .IN2(n1262), .Q(n1257) );
  AO21X1 U1111 ( .IN1(n989), .IN2(n1071), .IN3(n1264), .Q(n1262) );
  XOR2X1 U1112 ( .IN1(n1265), .IN2(n894), .Q(n1264) );
  NAND2X0 U1113 ( .IN1(n971), .IN2(n1079), .QN(n1265) );
  INVX0 U1114 ( .INP(n989), .ZN(n1079) );
  XOR2X1 U1115 ( .IN1(n1019), .IN2(n994), .Q(n1263) );
  NAND2X0 U1116 ( .IN1(n973), .IN2(n1022), .QN(n1255) );
  OA22X1 U1117 ( .IN1(n1106), .IN2(n1066), .IN3(n1063), .IN4(n1083), .Q(n1247)
         );
  INVX0 U1118 ( .INP(n1064), .ZN(n1083) );
  XNOR3X1 U1119 ( .IN1(n1266), .IN2(n1267), .IN3(n1004), .Q(n1066) );
  XOR3X1 U1120 ( .IN1(n1014), .IN2(n996), .IN3(n1009), .Q(n1267) );
  NOR2X0 U1121 ( .IN1(n1268), .IN2(n1269), .QN(n1266) );
  XOR2X1 U1122 ( .IN1(n1270), .IN2(n890), .Q(n1269) );
  NAND3X0 U1123 ( .IN1(n1022), .IN2(n1271), .IN3(n984), .QN(n1270) );
  AOI21X1 U1124 ( .IN1(n1022), .IN2(n984), .IN3(n1271), .QN(n1268) );
  XOR2X1 U1125 ( .IN1(n1253), .IN2(n1272), .Q(n1271) );
  XNOR3X1 U1126 ( .IN1(n1023), .IN2(n1273), .IN3(n1274), .Q(n1253) );
  XOR3X1 U1127 ( .IN1(n854), .IN2(n927), .IN3(n997), .Q(n1274) );
  XOR2X1 U1128 ( .IN1(n1017), .IN2(n993), .Q(n1273) );
  NOR2X0 U1129 ( .IN1(n1046), .IN2(n1064), .QN(n1106) );
  XNOR2X1 U1130 ( .IN1(n1275), .IN2(n1276), .Q(n1064) );
  OA22X1 U1131 ( .IN1(n1277), .IN2(n1278), .IN3(n1279), .IN4(n1280), .Q(n1276)
         );
  XNOR2X1 U1132 ( .IN1(n1281), .IN2(n1252), .Q(n1280) );
  AND2X1 U1133 ( .IN1(n1022), .IN2(n983), .Q(n1279) );
  NAND2X0 U1134 ( .IN1(n983), .IN2(n1022), .QN(n1278) );
  XOR2X1 U1135 ( .IN1(n1252), .IN2(n1281), .Q(n1277) );
  AO21X1 U1136 ( .IN1(n1282), .IN2(n1283), .IN3(n1284), .Q(n1252) );
  XOR2X1 U1137 ( .IN1(n963), .IN2(n1285), .Q(n1284) );
  NOR2X0 U1138 ( .IN1(n1283), .IN2(n1282), .QN(n1285) );
  XOR2X1 U1139 ( .IN1(n1176), .IN2(n1006), .Q(n1283) );
  INVX0 U1140 ( .INP(n978), .ZN(n1176) );
  XOR2X1 U1141 ( .IN1(n1029), .IN2(n1020), .Q(n1282) );
  INVX0 U1142 ( .INP(n979), .ZN(n1029) );
  OA21X1 U1143 ( .IN1(n1286), .IN2(n1287), .IN3(n1288), .Q(n1275) );
  XOR2X1 U1144 ( .IN1(n1289), .IN2(n893), .Q(n1288) );
  NAND2X0 U1145 ( .IN1(n1287), .IN2(n1286), .QN(n1289) );
  XOR2X1 U1146 ( .IN1(n1018), .IN2(n1002), .Q(n1287) );
  XOR2X1 U1147 ( .IN1(n1000), .IN2(n1012), .Q(n1286) );
  INVX0 U1148 ( .INP(n1063), .ZN(n1046) );
  XOR3X1 U1149 ( .IN1(n1290), .IN2(n1291), .IN3(n1292), .Q(n1063) );
  XOR2X1 U1150 ( .IN1(n1073), .IN2(n981), .Q(n1292) );
  INVX0 U1151 ( .INP(n980), .ZN(n1073) );
  OA21X1 U1152 ( .IN1(n1293), .IN2(n1294), .IN3(n1295), .Q(n1291) );
  NAND3X0 U1153 ( .IN1(n1022), .IN2(n1294), .IN3(n975), .QN(n1295) );
  XNOR2X1 U1154 ( .IN1(n1281), .IN2(n1272), .Q(n1294) );
  XOR3X1 U1155 ( .IN1(n1013), .IN2(n1296), .IN3(n1011), .Q(n1272) );
  OA21X1 U1156 ( .IN1(n1297), .IN2(n1056), .IN3(n1298), .Q(n1296) );
  XOR2X1 U1157 ( .IN1(n965), .IN2(n1299), .Q(n1298) );
  NOR2X0 U1158 ( .IN1(n1297), .IN2(n986), .QN(n1299) );
  INVX0 U1159 ( .INP(n972), .ZN(n1056) );
  XOR2X1 U1160 ( .IN1(n1300), .IN2(n895), .Q(n1297) );
  NAND2X0 U1161 ( .IN1(n972), .IN2(n987), .QN(n1300) );
  AO21X1 U1162 ( .IN1(n1301), .IN2(n1302), .IN3(n1303), .Q(n1281) );
  XOR2X1 U1163 ( .IN1(n1304), .IN2(n892), .Q(n1303) );
  OR2X1 U1164 ( .IN1(n1302), .IN2(n1301), .Q(n1304) );
  XOR2X1 U1165 ( .IN1(n1015), .IN2(n991), .Q(n1302) );
  XOR2X1 U1166 ( .IN1(n1016), .IN2(n1133), .Q(n1301) );
  INVX0 U1167 ( .INP(n1003), .ZN(n1133) );
  NOR2X0 U1168 ( .IN1(n1021), .IN2(n974), .QN(n1293) );
  OA21X1 U1169 ( .IN1(n988), .IN2(n1007), .IN3(n1305), .Q(n1290) );
  XOR2X1 U1170 ( .IN1(n964), .IN2(n1306), .Q(n1305) );
  NOR2X0 U1171 ( .IN1(n1008), .IN2(n1134), .QN(n1306) );
  INVX0 U1172 ( .INP(n1052), .ZN(n1040) );
  XOR3X1 U1173 ( .IN1(n1307), .IN2(n1308), .IN3(n986), .Q(n1052) );
  XOR3X1 U1174 ( .IN1(n978), .IN2(n1017), .IN3(n991), .Q(n1308) );
  OA22X1 U1175 ( .IN1(n1309), .IN2(n1310), .IN3(n1311), .IN4(n1312), .Q(n1307)
         );
  XNOR2X1 U1176 ( .IN1(n1313), .IN2(n1314), .Q(n1312) );
  AND2X1 U1177 ( .IN1(n1022), .IN2(n982), .Q(n1311) );
  NAND2X0 U1178 ( .IN1(n982), .IN2(n1022), .QN(n1310) );
  XOR2X1 U1179 ( .IN1(n1314), .IN2(n1313), .Q(n1309) );
  AO21X1 U1180 ( .IN1(n1315), .IN2(n1316), .IN3(n1317), .Q(n1044) );
  XOR3X1 U1181 ( .IN1(n1318), .IN2(n1319), .IN3(n1320), .Q(n1317) );
  XOR2X1 U1182 ( .IN1(n1246), .IN2(n1314), .Q(n1320) );
  AOI21X1 U1183 ( .IN1(n1321), .IN2(n1322), .IN3(n1323), .QN(n1314) );
  XOR2X1 U1184 ( .IN1(n962), .IN2(n1324), .Q(n1323) );
  NOR2X0 U1185 ( .IN1(n1321), .IN2(n1322), .QN(n1324) );
  AO21X1 U1186 ( .IN1(n1002), .IN2(n995), .IN3(n1325), .Q(n1322) );
  XOR2X1 U1187 ( .IN1(n966), .IN2(n1326), .Q(n1325) );
  NOR2X0 U1188 ( .IN1(n1002), .IN2(n995), .QN(n1326) );
  XOR2X1 U1189 ( .IN1(n1134), .IN2(n994), .Q(n1321) );
  INVX0 U1190 ( .INP(n988), .ZN(n1134) );
  XOR3X1 U1191 ( .IN1(n1019), .IN2(n1008), .IN3(n1327), .Q(n1246) );
  XNOR2X1 U1192 ( .IN1(n1014), .IN2(n1018), .Q(n1327) );
  NOR2X0 U1193 ( .IN1(n1315), .IN2(n1316), .QN(n1319) );
  AND2X1 U1194 ( .IN1(n970), .IN2(n1022), .Q(n1318) );
  INVX0 U1195 ( .INP(n814), .ZN(n1316) );
  AOI21X1 U1196 ( .IN1(n1328), .IN2(n1329), .IN3(n1330), .QN(n1315) );
  XOR2X1 U1197 ( .IN1(n1331), .IN2(n891), .Q(n1330) );
  NAND2X0 U1198 ( .IN1(n1332), .IN2(n1333), .QN(n1331) );
  XOR2X1 U1199 ( .IN1(n1003), .IN2(n1011), .Q(n1333) );
  XOR2X1 U1200 ( .IN1(n1023), .IN2(n1162), .Q(n1332) );
  INVX0 U1201 ( .INP(n1020), .ZN(n1162) );
  XOR2X1 U1202 ( .IN1(n1020), .IN2(n1023), .Q(n1329) );
  XOR2X1 U1203 ( .IN1(n1010), .IN2(n1003), .Q(n1328) );
  XOR2X1 U1204 ( .IN1(n1334), .IN2(n1335), .Q(n1031) );
  XOR3X1 U1205 ( .IN1(n1016), .IN2(n1013), .IN3(n1336), .Q(n1335) );
  OA21X1 U1206 ( .IN1(n1337), .IN2(n1338), .IN3(n1339), .Q(n1336) );
  NAND3X0 U1207 ( .IN1(n1022), .IN2(n1338), .IN3(n977), .QN(n1339) );
  XOR2X1 U1208 ( .IN1(n1245), .IN2(n1313), .Q(n1338) );
  XNOR3X1 U1209 ( .IN1(n1004), .IN2(n989), .IN3(n1340), .Q(n1313) );
  XOR2X1 U1210 ( .IN1(n1161), .IN2(n1012), .Q(n1340) );
  INVX0 U1211 ( .INP(n981), .ZN(n1161) );
  XOR3X1 U1212 ( .IN1(n1071), .IN2(n980), .IN3(n1341), .Q(n1245) );
  XOR3X1 U1213 ( .IN1(n855), .IN2(n999), .IN3(n1009), .Q(n1341) );
  INVX0 U1214 ( .INP(n971), .ZN(n1071) );
  NOR2X0 U1215 ( .IN1(n1021), .IN2(n976), .QN(n1337) );
  XOR3X1 U1216 ( .IN1(n853), .IN2(n979), .IN3(n992), .Q(n1334) );
endmodule

