
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762;

  XNOR2X1 U415 ( .IN1(n390), .IN2(keyinput126), .Q(G1342) );
  NAND2X0 U416 ( .IN1(n391), .IN2(n392), .QN(n390) );
  NAND3X0 U417 ( .IN1(n393), .IN2(n394), .IN3(n395), .QN(n392) );
  XOR2X1 U418 ( .IN1(n396), .IN2(keyinput103), .Q(n391) );
  NAND2X0 U419 ( .IN1(G19), .IN2(n394), .QN(n396) );
  XNOR2X1 U420 ( .IN1(n397), .IN2(keyinput94), .Q(n394) );
  NAND3X0 U421 ( .IN1(n393), .IN2(G19), .IN3(n395), .QN(n397) );
  XOR2X1 U422 ( .IN1(n398), .IN2(G32), .Q(G1355) );
  NAND2X0 U423 ( .IN1(n399), .IN2(n400), .QN(n398) );
  OA21X1 U424 ( .IN1(n401), .IN2(n402), .IN3(n403), .Q(G1354) );
  XOR2X1 U425 ( .IN1(keyinput112), .IN2(n404), .Q(n403) );
  NOR2X0 U426 ( .IN1(n402), .IN2(n405), .QN(n404) );
  XOR2X1 U427 ( .IN1(n406), .IN2(keyinput96), .Q(n402) );
  OR2X1 U428 ( .IN1(n405), .IN2(n401), .Q(n406) );
  XOR2X1 U429 ( .IN1(n407), .IN2(keyinput91), .Q(n401) );
  NAND2X0 U430 ( .IN1(n399), .IN2(n393), .QN(n407) );
  OA21X1 U431 ( .IN1(n408), .IN2(n409), .IN3(n410), .Q(G1353) );
  XOR2X1 U432 ( .IN1(n411), .IN2(keyinput111), .Q(n410) );
  NAND2X0 U433 ( .IN1(n408), .IN2(n409), .QN(n411) );
  XOR2X1 U434 ( .IN1(n412), .IN2(keyinput90), .Q(n408) );
  NAND2X0 U435 ( .IN1(n399), .IN2(n413), .QN(n412) );
  OA21X1 U436 ( .IN1(n414), .IN2(n415), .IN3(n416), .Q(G1350) );
  XOR2X1 U437 ( .IN1(keyinput109), .IN2(n417), .Q(n416) );
  AND2X1 U438 ( .IN1(n414), .IN2(n415), .Q(n417) );
  XNOR2X1 U439 ( .IN1(n418), .IN2(keyinput88), .Q(n415) );
  NAND2X0 U440 ( .IN1(n419), .IN2(n393), .QN(n418) );
  OA21X1 U441 ( .IN1(n420), .IN2(n421), .IN3(n422), .Q(G1349) );
  XOR2X1 U442 ( .IN1(n423), .IN2(keyinput108), .Q(n422) );
  NAND2X0 U443 ( .IN1(n420), .IN2(n421), .QN(n423) );
  XOR2X1 U444 ( .IN1(n424), .IN2(keyinput87), .Q(n420) );
  NAND2X0 U445 ( .IN1(n419), .IN2(n413), .QN(n424) );
  OA21X1 U446 ( .IN1(n425), .IN2(n426), .IN3(n427), .Q(G1348) );
  XOR2X1 U447 ( .IN1(n428), .IN2(keyinput107), .Q(n427) );
  NAND2X0 U448 ( .IN1(G25), .IN2(n429), .QN(n428) );
  INVX0 U449 ( .INP(n425), .ZN(n429) );
  INVX0 U450 ( .INP(n430), .ZN(n426) );
  XOR2X1 U451 ( .IN1(n431), .IN2(keyinput95), .Q(n425) );
  NAND2X0 U452 ( .IN1(n430), .IN2(G25), .QN(n431) );
  XOR2X1 U453 ( .IN1(n432), .IN2(keyinput86), .Q(n430) );
  NAND2X0 U454 ( .IN1(n419), .IN2(n433), .QN(n432) );
  NOR2X0 U455 ( .IN1(n434), .IN2(n435), .QN(G1347) );
  XOR2X1 U456 ( .IN1(keyinput106), .IN2(n436), .Q(n435) );
  NOR2X0 U457 ( .IN1(n437), .IN2(n438), .QN(n436) );
  NOR3X0 U458 ( .IN1(n439), .IN2(n437), .IN3(n440), .QN(n434) );
  NOR3X0 U459 ( .IN1(n440), .IN2(n438), .IN3(n439), .QN(n437) );
  INVX0 U460 ( .INP(G24), .ZN(n438) );
  NOR2X0 U461 ( .IN1(n441), .IN2(n442), .QN(G1344) );
  XOR2X1 U462 ( .IN1(keyinput104), .IN2(n443), .Q(n442) );
  NOR2X0 U463 ( .IN1(n444), .IN2(n445), .QN(n443) );
  NOR3X0 U464 ( .IN1(n439), .IN2(n444), .IN3(n446), .QN(n441) );
  NOR3X0 U465 ( .IN1(n445), .IN2(n446), .IN3(n439), .QN(n444) );
  XOR3X1 U466 ( .IN1(keyinput84), .IN2(G18), .IN3(n447), .Q(G1341) );
  NAND2X0 U467 ( .IN1(n395), .IN2(n413), .QN(n447) );
  XOR3X1 U468 ( .IN1(keyinput82), .IN2(G16), .IN3(n448), .Q(G1339) );
  NOR2X0 U469 ( .IN1(n449), .IN2(n450), .QN(n448) );
  NOR2X0 U470 ( .IN1(n451), .IN2(n452), .QN(G1337) );
  XOR2X1 U471 ( .IN1(n453), .IN2(keyinput102), .Q(n452) );
  NAND3X0 U472 ( .IN1(n454), .IN2(n455), .IN3(n456), .QN(n453) );
  OA21X1 U473 ( .IN1(n457), .IN2(n450), .IN3(G14), .Q(n451) );
  OA22X1 U474 ( .IN1(n458), .IN2(n459), .IN3(n458), .IN4(n460), .Q(G1334) );
  XOR2X1 U475 ( .IN1(n461), .IN2(keyinput93), .Q(n458) );
  OR2X1 U476 ( .IN1(n459), .IN2(n460), .Q(n461) );
  NAND2X0 U477 ( .IN1(n462), .IN2(n463), .QN(n459) );
  XOR3X1 U478 ( .IN1(keyinput80), .IN2(G10), .IN3(n464), .Q(G1333) );
  NOR2X0 U479 ( .IN1(n457), .IN2(n465), .QN(n464) );
  OA22X1 U480 ( .IN1(n466), .IN2(n467), .IN3(n468), .IN4(n467), .Q(G1332) );
  XNOR2X1 U481 ( .IN1(n469), .IN2(keyinput92), .Q(n467) );
  OR2X1 U482 ( .IN1(n466), .IN2(n468), .Q(n469) );
  NAND2X0 U483 ( .IN1(n463), .IN2(n470), .QN(n466) );
  OA21X1 U484 ( .IN1(G7), .IN2(n471), .IN3(n472), .Q(G1330) );
  XOR2X1 U485 ( .IN1(keyinput99), .IN2(n473), .Q(n472) );
  NOR2X0 U486 ( .IN1(n474), .IN2(n475), .QN(n473) );
  INVX0 U487 ( .INP(n474), .ZN(n471) );
  NOR2X0 U488 ( .IN1(n476), .IN2(n477), .QN(n474) );
  XOR2X1 U489 ( .IN1(keyinput115), .IN2(n478), .Q(G1329) );
  MUX21X1 U490 ( .IN1(n479), .IN2(n480), .S(G6), .Q(n478) );
  OR2X1 U491 ( .IN1(n476), .IN2(n457), .Q(n480) );
  NOR2X0 U492 ( .IN1(n457), .IN2(n476), .QN(n479) );
  XOR2X1 U493 ( .IN1(n481), .IN2(n482), .Q(G1328) );
  NOR2X0 U494 ( .IN1(n483), .IN2(n476), .QN(n482) );
  XNOR2X1 U495 ( .IN1(keyinput114), .IN2(n484), .Q(G1327) );
  OA21X1 U496 ( .IN1(keyinput98), .IN2(G4), .IN3(n485), .Q(n484) );
  XOR2X1 U497 ( .IN1(n486), .IN2(n487), .Q(n485) );
  NOR2X0 U498 ( .IN1(n449), .IN2(n488), .QN(n487) );
  NAND2X0 U499 ( .IN1(keyinput98), .IN2(G4), .QN(n486) );
  XNOR2X1 U500 ( .IN1(G2), .IN2(n489), .Q(G1325) );
  NOR2X0 U501 ( .IN1(n457), .IN2(n488), .QN(n489) );
  XOR3X1 U502 ( .IN1(keyinput79), .IN2(G1), .IN3(n490), .Q(G1324) );
  NAND2X0 U503 ( .IN1(n491), .IN2(n470), .QN(n490) );
  XOR2X1 U504 ( .IN1(keyinput120), .IN2(n492), .Q(G1345) );
  MUX21X1 U505 ( .IN1(n493), .IN2(n494), .S(G22), .Q(n492) );
  NAND2X0 U506 ( .IN1(n495), .IN2(n413), .QN(n494) );
  NOR2X0 U507 ( .IN1(n496), .IN2(n439), .QN(n493) );
  XOR2X1 U508 ( .IN1(keyinput119), .IN2(n497), .Q(G1343) );
  MUX21X1 U509 ( .IN1(n498), .IN2(n499), .S(G20), .Q(n497) );
  NAND2X0 U510 ( .IN1(n395), .IN2(n400), .QN(n499) );
  NOR2X0 U511 ( .IN1(n440), .IN2(n500), .QN(n498) );
  XOR2X1 U512 ( .IN1(keyinput116), .IN2(n501), .Q(G1335) );
  MUX21X1 U513 ( .IN1(n502), .IN2(n503), .S(G12), .Q(n501) );
  NAND2X0 U514 ( .IN1(n463), .IN2(n504), .QN(n503) );
  INVX0 U515 ( .INP(n465), .ZN(n463) );
  NOR2X0 U516 ( .IN1(n449), .IN2(n465), .QN(n502) );
  XOR2X1 U517 ( .IN1(n505), .IN2(keyinput78), .Q(n465) );
  NAND3X0 U518 ( .IN1(n446), .IN2(n413), .IN3(n506), .QN(n505) );
  XOR2X1 U519 ( .IN1(keyinput122), .IN2(n507), .Q(G1352) );
  OA21X1 U520 ( .IN1(n508), .IN2(n509), .IN3(n510), .Q(n507) );
  XOR2X1 U521 ( .IN1(n511), .IN2(keyinput110), .Q(n510) );
  NAND3X0 U522 ( .IN1(n433), .IN2(n509), .IN3(n399), .QN(n511) );
  INVX0 U523 ( .INP(n512), .ZN(n399) );
  INVX0 U524 ( .INP(G29), .ZN(n509) );
  NOR2X0 U525 ( .IN1(n446), .IN2(n512), .QN(n508) );
  NAND3X0 U526 ( .IN1(n513), .IN2(n454), .IN3(n483), .QN(n512) );
  XOR3X1 U527 ( .IN1(n514), .IN2(n515), .IN3(n516), .Q(G1351) );
  NAND2X0 U528 ( .IN1(n419), .IN2(n400), .QN(n516) );
  AND4X1 U529 ( .IN1(n454), .IN2(n517), .IN3(n462), .IN4(n518), .Q(n419) );
  NOR2X0 U530 ( .IN1(n504), .IN2(n519), .QN(n518) );
  XOR2X1 U531 ( .IN1(keyinput76), .IN2(n483), .Q(n519) );
  XOR2X1 U532 ( .IN1(keyinput89), .IN2(keyinput127), .Q(n514) );
  XOR2X1 U533 ( .IN1(keyinput121), .IN2(n520), .Q(G1346) );
  OA21X1 U534 ( .IN1(n521), .IN2(n522), .IN3(n523), .Q(n520) );
  XOR2X1 U535 ( .IN1(n524), .IN2(keyinput105), .Q(n523) );
  NAND2X0 U536 ( .IN1(n521), .IN2(n522), .QN(n524) );
  INVX0 U537 ( .INP(G23), .ZN(n522) );
  XOR2X1 U538 ( .IN1(n525), .IN2(keyinput85), .Q(n521) );
  NAND2X0 U539 ( .IN1(n495), .IN2(n393), .QN(n525) );
  INVX0 U540 ( .INP(n439), .ZN(n495) );
  NAND3X0 U541 ( .IN1(n457), .IN2(n470), .IN3(n513), .QN(n439) );
  AND3X1 U542 ( .IN1(n517), .IN2(n504), .IN3(n477), .Q(n513) );
  XNOR3X1 U543 ( .IN1(n526), .IN2(G17), .IN3(n527), .Q(G1340) );
  NAND2X0 U544 ( .IN1(n395), .IN2(n433), .QN(n527) );
  INVX0 U545 ( .INP(n500), .ZN(n395) );
  NAND4X0 U546 ( .IN1(n517), .IN2(n470), .IN3(n528), .IN4(n529), .QN(n500) );
  NOR2X0 U547 ( .IN1(n504), .IN2(n477), .QN(n529) );
  XOR2X1 U548 ( .IN1(keyinput75), .IN2(n454), .Q(n528) );
  NAND2X0 U549 ( .IN1(n530), .IN2(n531), .QN(n517) );
  NAND3X0 U550 ( .IN1(n532), .IN2(n446), .IN3(n533), .QN(n531) );
  XOR2X1 U551 ( .IN1(n534), .IN2(n440), .Q(n533) );
  NAND2X0 U552 ( .IN1(keyinput73), .IN2(n413), .QN(n534) );
  NAND3X0 U553 ( .IN1(n496), .IN2(n440), .IN3(n535), .QN(n530) );
  XOR2X1 U554 ( .IN1(n393), .IN2(n536), .Q(n535) );
  NOR2X0 U555 ( .IN1(keyinput74), .IN2(n446), .QN(n536) );
  XOR2X1 U556 ( .IN1(keyinput83), .IN2(keyinput125), .Q(n526) );
  XOR2X1 U557 ( .IN1(n537), .IN2(keyinput118), .Q(G1338) );
  MUX21X1 U558 ( .IN1(n538), .IN2(n539), .S(G15), .Q(n537) );
  NOR2X0 U559 ( .IN1(n477), .IN2(n450), .QN(n539) );
  NAND2X0 U560 ( .IN1(n456), .IN2(n462), .QN(n538) );
  XOR3X1 U561 ( .IN1(keyinput124), .IN2(keyinput117), .IN3(n540), .Q(G1336) );
  OA21X1 U562 ( .IN1(n541), .IN2(n542), .IN3(n543), .Q(n540) );
  XOR2X1 U563 ( .IN1(n544), .IN2(keyinput101), .Q(n543) );
  NAND2X0 U564 ( .IN1(n541), .IN2(n542), .QN(n544) );
  XOR2X1 U565 ( .IN1(n545), .IN2(keyinput81), .Q(n541) );
  NAND2X0 U566 ( .IN1(n456), .IN2(n470), .QN(n545) );
  INVX0 U567 ( .INP(n450), .ZN(n456) );
  NAND4X0 U568 ( .IN1(n413), .IN2(n546), .IN3(n400), .IN4(n547), .QN(n450) );
  NOR2X0 U569 ( .IN1(n433), .IN2(n548), .QN(n547) );
  XOR2X1 U570 ( .IN1(keyinput72), .IN2(n532), .Q(n548) );
  XOR2X1 U571 ( .IN1(keyinput123), .IN2(n549), .Q(G1331) );
  OA21X1 U572 ( .IN1(keyinput100), .IN2(G8), .IN3(n550), .Q(n549) );
  XOR2X1 U573 ( .IN1(n551), .IN2(n552), .Q(n550) );
  NOR2X0 U574 ( .IN1(n449), .IN2(n476), .QN(n552) );
  NAND4X0 U575 ( .IN1(n400), .IN2(n496), .IN3(n553), .IN4(n433), .QN(n476) );
  AND2X1 U576 ( .IN1(n546), .IN2(n532), .Q(n553) );
  INVX0 U577 ( .INP(n393), .ZN(n532) );
  NAND2X0 U578 ( .IN1(keyinput100), .IN2(G8), .QN(n551) );
  XOR2X1 U579 ( .IN1(keyinput113), .IN2(n554), .Q(G1326) );
  OA21X1 U580 ( .IN1(n555), .IN2(n556), .IN3(n557), .Q(n554) );
  XOR2X1 U581 ( .IN1(n558), .IN2(keyinput97), .Q(n557) );
  NAND3X0 U582 ( .IN1(n491), .IN2(n556), .IN3(n462), .QN(n558) );
  INVX0 U583 ( .INP(n488), .ZN(n491) );
  NOR2X0 U584 ( .IN1(n488), .IN2(n477), .QN(n555) );
  XOR2X1 U585 ( .IN1(n559), .IN2(keyinput77), .Q(n488) );
  NAND3X0 U586 ( .IN1(n560), .IN2(n433), .IN3(n506), .QN(n559) );
  AND3X1 U587 ( .IN1(n440), .IN2(n546), .IN3(n393), .Q(n506) );
  XOR3X1 U588 ( .IN1(keyinput69), .IN2(n561), .IN3(n562), .Q(n393) );
  MUX21X1 U589 ( .IN1(n563), .IN2(n564), .S(n565), .Q(n562) );
  OA21X1 U590 ( .IN1(n566), .IN2(n567), .IN3(n568), .Q(n565) );
  XOR2X1 U591 ( .IN1(n569), .IN2(keyinput48), .Q(n568) );
  NAND2X0 U592 ( .IN1(n566), .IN2(n567), .QN(n569) );
  AND2X1 U593 ( .IN1(G41), .IN2(G39), .Q(n564) );
  NAND2X0 U594 ( .IN1(G39), .IN2(G41), .QN(n563) );
  OA21X1 U595 ( .IN1(n570), .IN2(n571), .IN3(n572), .Q(n561) );
  XOR2X1 U596 ( .IN1(n573), .IN2(keyinput43), .Q(n572) );
  NAND2X0 U597 ( .IN1(n570), .IN2(n571), .QN(n573) );
  XOR3X1 U598 ( .IN1(keyinput33), .IN2(G23), .IN3(G19), .Q(n571) );
  XOR2X1 U599 ( .IN1(n405), .IN2(G27), .Q(n570) );
  NAND2X0 U600 ( .IN1(n574), .IN2(n575), .QN(n546) );
  NAND3X0 U601 ( .IN1(n457), .IN2(n576), .IN3(n483), .QN(n575) );
  NAND2X0 U602 ( .IN1(n462), .IN2(n504), .QN(n576) );
  NAND3X0 U603 ( .IN1(n449), .IN2(n477), .IN3(n577), .QN(n574) );
  XOR2X1 U604 ( .IN1(n578), .IN2(n483), .Q(n577) );
  INVX0 U605 ( .INP(n470), .ZN(n483) );
  AO22X1 U606 ( .IN1(n579), .IN2(n580), .IN3(n581), .IN4(n582), .Q(n470) );
  INVX0 U607 ( .INP(keyinput63), .ZN(n582) );
  NAND2X0 U608 ( .IN1(n583), .IN2(n580), .QN(n581) );
  NAND2X0 U609 ( .IN1(n584), .IN2(n583), .QN(n580) );
  AO21X1 U610 ( .IN1(keyinput63), .IN2(n583), .IN3(n584), .Q(n579) );
  XOR2X1 U611 ( .IN1(n585), .IN2(keyinput58), .Q(n584) );
  OAI21X1 U612 ( .IN1(n586), .IN2(n587), .IN3(n588), .QN(n585) );
  XNOR2X1 U613 ( .IN1(n589), .IN2(keyinput53), .Q(n588) );
  NAND2X0 U614 ( .IN1(n587), .IN2(n586), .QN(n589) );
  XNOR2X1 U615 ( .IN1(n590), .IN2(keyinput0), .Q(n587) );
  NAND2X0 U616 ( .IN1(G33), .IN2(G41), .QN(n590) );
  AO21X1 U617 ( .IN1(n591), .IN2(n592), .IN3(n593), .Q(n586) );
  XOR2X1 U618 ( .IN1(n594), .IN2(keyinput50), .Q(n593) );
  OR2X1 U619 ( .IN1(n591), .IN2(n592), .Q(n594) );
  INVX0 U620 ( .INP(n595), .ZN(n591) );
  AO21X1 U621 ( .IN1(n596), .IN2(n597), .IN3(n598), .Q(n583) );
  XOR2X1 U622 ( .IN1(keyinput40), .IN2(n599), .Q(n598) );
  NOR2X0 U623 ( .IN1(n596), .IN2(n597), .QN(n599) );
  AO21X1 U624 ( .IN1(G13), .IN2(n468), .IN3(n600), .Q(n597) );
  XOR2X1 U625 ( .IN1(n601), .IN2(keyinput21), .Q(n600) );
  NAND2X0 U626 ( .IN1(G9), .IN2(n542), .QN(n601) );
  INVX0 U627 ( .INP(G13), .ZN(n542) );
  AOI21X1 U628 ( .IN1(n602), .IN2(G1), .IN3(n603), .QN(n596) );
  XOR2X1 U629 ( .IN1(n604), .IN2(keyinput20), .Q(n603) );
  NAND2X0 U630 ( .IN1(n602), .IN2(G5), .QN(n604) );
  XOR2X1 U631 ( .IN1(n605), .IN2(keyinput9), .Q(n602) );
  NAND2X0 U632 ( .IN1(G5), .IN2(G1), .QN(n605) );
  NAND2X0 U633 ( .IN1(keyinput70), .IN2(n454), .QN(n578) );
  INVX0 U634 ( .INP(n457), .ZN(n454) );
  XOR3X1 U635 ( .IN1(n606), .IN2(n607), .IN3(n608), .Q(n457) );
  NAND2X0 U636 ( .IN1(n609), .IN2(n610), .QN(n608) );
  XOR2X1 U637 ( .IN1(n611), .IN2(keyinput56), .Q(n610) );
  NAND2X0 U638 ( .IN1(n612), .IN2(n613), .QN(n611) );
  XOR2X1 U639 ( .IN1(n614), .IN2(n615), .Q(n613) );
  XOR2X1 U640 ( .IN1(n616), .IN2(keyinput1), .Q(n612) );
  XOR2X1 U641 ( .IN1(n617), .IN2(keyinput55), .Q(n609) );
  NAND2X0 U642 ( .IN1(n618), .IN2(n619), .QN(n617) );
  XNOR2X1 U643 ( .IN1(keyinput1), .IN2(n616), .Q(n619) );
  NAND2X0 U644 ( .IN1(G34), .IN2(G41), .QN(n616) );
  XOR2X1 U645 ( .IN1(n620), .IN2(n615), .Q(n618) );
  XOR2X1 U646 ( .IN1(G6), .IN2(G2), .Q(n607) );
  OA21X1 U647 ( .IN1(G10), .IN2(n455), .IN3(n621), .Q(n606) );
  XOR2X1 U648 ( .IN1(n622), .IN2(keyinput22), .Q(n621) );
  NAND2X0 U649 ( .IN1(G10), .IN2(n455), .QN(n622) );
  INVX0 U650 ( .INP(G14), .ZN(n455) );
  INVX0 U651 ( .INP(n462), .ZN(n477) );
  XNOR2X1 U652 ( .IN1(keyinput67), .IN2(n623), .Q(n462) );
  OA21X1 U653 ( .IN1(n624), .IN2(n625), .IN3(n626), .Q(n623) );
  XOR2X1 U654 ( .IN1(keyinput64), .IN2(n627), .Q(n626) );
  AND2X1 U655 ( .IN1(n625), .IN2(n624), .Q(n627) );
  XNOR3X1 U656 ( .IN1(keyinput59), .IN2(keyinput2), .IN3(n628), .Q(n625) );
  XOR2X1 U657 ( .IN1(n629), .IN2(n630), .Q(n628) );
  OA21X1 U658 ( .IN1(n595), .IN2(n615), .IN3(n631), .Q(n630) );
  XOR2X1 U659 ( .IN1(keyinput51), .IN2(n632), .Q(n631) );
  AND2X1 U660 ( .IN1(n615), .IN2(n595), .Q(n632) );
  XOR3X1 U661 ( .IN1(G26), .IN2(n633), .IN3(G25), .Q(n615) );
  OA21X1 U662 ( .IN1(G27), .IN2(G28), .IN3(n634), .Q(n633) );
  XOR2X1 U663 ( .IN1(keyinput8), .IN2(n635), .Q(n634) );
  NOR2X0 U664 ( .IN1(n515), .IN2(n414), .QN(n635) );
  INVX0 U665 ( .INP(G27), .ZN(n414) );
  XNOR3X1 U666 ( .IN1(keyinput30), .IN2(n636), .IN3(n637), .Q(n595) );
  OA21X1 U667 ( .IN1(G19), .IN2(G20), .IN3(n638), .Q(n637) );
  XOR2X1 U668 ( .IN1(keyinput7), .IN2(n639), .Q(n638) );
  AND2X1 U669 ( .IN1(G19), .IN2(G20), .Q(n639) );
  OA21X1 U670 ( .IN1(G17), .IN2(n640), .IN3(n641), .Q(n636) );
  XOR2X1 U671 ( .IN1(keyinput18), .IN2(n642), .Q(n641) );
  AND2X1 U672 ( .IN1(n640), .IN2(G17), .Q(n642) );
  NAND2X0 U673 ( .IN1(G35), .IN2(G41), .QN(n629) );
  OA21X1 U674 ( .IN1(n643), .IN2(n644), .IN3(n645), .Q(n624) );
  XOR2X1 U675 ( .IN1(n646), .IN2(keyinput41), .Q(n645) );
  NAND3X0 U676 ( .IN1(n647), .IN2(n648), .IN3(n644), .QN(n646) );
  NAND2X0 U677 ( .IN1(G3), .IN2(n475), .QN(n648) );
  XNOR2X1 U678 ( .IN1(keyinput31), .IN2(n649), .Q(n644) );
  OA21X1 U679 ( .IN1(G15), .IN2(G11), .IN3(n650), .Q(n649) );
  XOR2X1 U680 ( .IN1(keyinput10), .IN2(n651), .Q(n650) );
  NOR2X0 U681 ( .IN1(n652), .IN2(n460), .QN(n651) );
  INVX0 U682 ( .INP(G11), .ZN(n460) );
  OA21X1 U683 ( .IN1(G7), .IN2(n556), .IN3(n647), .Q(n643) );
  XOR2X1 U684 ( .IN1(n653), .IN2(keyinput23), .Q(n647) );
  NAND2X0 U685 ( .IN1(G7), .IN2(n556), .QN(n653) );
  INVX0 U686 ( .INP(n504), .ZN(n449) );
  NAND2X0 U687 ( .IN1(n654), .IN2(n655), .QN(n504) );
  NAND3X0 U688 ( .IN1(n656), .IN2(n657), .IN3(n658), .QN(n655) );
  XOR2X1 U689 ( .IN1(keyinput65), .IN2(n659), .Q(n654) );
  AND2X1 U690 ( .IN1(n656), .IN2(n660), .Q(n659) );
  NAND3X0 U691 ( .IN1(n660), .IN2(n657), .IN3(n658), .QN(n656) );
  XOR2X1 U692 ( .IN1(n661), .IN2(keyinput54), .Q(n658) );
  NAND3X0 U693 ( .IN1(G41), .IN2(G36), .IN3(n662), .QN(n661) );
  AO21X1 U694 ( .IN1(G41), .IN2(G36), .IN3(n662), .Q(n657) );
  XOR2X1 U695 ( .IN1(n620), .IN2(n592), .Q(n662) );
  XOR3X1 U696 ( .IN1(G24), .IN2(n663), .IN3(G23), .Q(n592) );
  OA21X1 U697 ( .IN1(G22), .IN2(n445), .IN3(n664), .Q(n663) );
  XOR2X1 U698 ( .IN1(keyinput19), .IN2(n665), .Q(n664) );
  NOR2X0 U699 ( .IN1(G21), .IN2(n666), .QN(n665) );
  INVX0 U700 ( .INP(G22), .ZN(n666) );
  INVX0 U701 ( .INP(n614), .ZN(n620) );
  XNOR3X1 U702 ( .IN1(G30), .IN2(G29), .IN3(n667), .Q(n614) );
  XOR2X1 U703 ( .IN1(G32), .IN2(n405), .Q(n667) );
  INVX0 U704 ( .INP(G31), .ZN(n405) );
  XNOR3X1 U705 ( .IN1(keyinput32), .IN2(G8), .IN3(n668), .Q(n660) );
  XNOR2X1 U706 ( .IN1(G4), .IN2(n669), .Q(n668) );
  OA21X1 U707 ( .IN1(G16), .IN2(G12), .IN3(n670), .Q(n669) );
  XOR2X1 U708 ( .IN1(keyinput11), .IN2(n671), .Q(n670) );
  NOR2X0 U709 ( .IN1(n672), .IN2(n673), .QN(n671) );
  INVX0 U710 ( .INP(n400), .ZN(n440) );
  XNOR2X1 U711 ( .IN1(keyinput68), .IN2(n674), .Q(n400) );
  OA21X1 U712 ( .IN1(n675), .IN2(n676), .IN3(n677), .Q(n674) );
  XOR2X1 U713 ( .IN1(n678), .IN2(keyinput62), .Q(n677) );
  NAND2X0 U714 ( .IN1(n675), .IN2(n676), .QN(n678) );
  AO21X1 U715 ( .IN1(n679), .IN2(n680), .IN3(n681), .Q(n676) );
  XOR2X1 U716 ( .IN1(keyinput57), .IN2(n682), .Q(n681) );
  NOR2X0 U717 ( .IN1(n679), .IN2(n680), .QN(n682) );
  AO21X1 U718 ( .IN1(n683), .IN2(n684), .IN3(n685), .Q(n680) );
  XOR2X1 U719 ( .IN1(keyinput49), .IN2(n686), .Q(n685) );
  AND2X1 U720 ( .IN1(n687), .IN2(n683), .Q(n686) );
  XNOR2X1 U721 ( .IN1(n688), .IN2(keyinput47), .Q(n683) );
  NAND2X0 U722 ( .IN1(n687), .IN2(n684), .QN(n688) );
  NAND2X0 U723 ( .IN1(G40), .IN2(G41), .QN(n679) );
  XNOR3X1 U724 ( .IN1(keyinput34), .IN2(G32), .IN3(n689), .Q(n675) );
  XOR2X1 U725 ( .IN1(n515), .IN2(n690), .Q(n689) );
  OA21X1 U726 ( .IN1(G24), .IN2(G20), .IN3(n691), .Q(n690) );
  XOR2X1 U727 ( .IN1(n692), .IN2(keyinput12), .Q(n691) );
  NAND2X0 U728 ( .IN1(G20), .IN2(G24), .QN(n692) );
  INVX0 U729 ( .INP(G28), .ZN(n515) );
  INVX0 U730 ( .INP(n446), .ZN(n433) );
  XOR2X1 U731 ( .IN1(n693), .IN2(n694), .Q(n446) );
  XNOR3X1 U732 ( .IN1(n695), .IN2(n696), .IN3(n697), .Q(n694) );
  NAND2X0 U733 ( .IN1(G37), .IN2(G41), .QN(n697) );
  OA21X1 U734 ( .IN1(n698), .IN2(n699), .IN3(n700), .Q(n696) );
  XOR2X1 U735 ( .IN1(keyinput35), .IN2(n701), .Q(n700) );
  AND2X1 U736 ( .IN1(n699), .IN2(n698), .Q(n701) );
  NAND2X0 U737 ( .IN1(n702), .IN2(n703), .QN(n699) );
  XOR2X1 U738 ( .IN1(keyinput25), .IN2(n704), .Q(n703) );
  NOR2X0 U739 ( .IN1(G17), .IN2(n445), .QN(n704) );
  XOR2X1 U740 ( .IN1(n705), .IN2(keyinput24), .Q(n702) );
  NAND2X0 U741 ( .IN1(G17), .IN2(n445), .QN(n705) );
  INVX0 U742 ( .INP(G21), .ZN(n445) );
  XOR2X1 U743 ( .IN1(G25), .IN2(G29), .Q(n698) );
  OA21X1 U744 ( .IN1(n706), .IN2(n684), .IN3(n707), .Q(n695) );
  XOR2X1 U745 ( .IN1(keyinput46), .IN2(n708), .Q(n707) );
  NOR2X0 U746 ( .IN1(n566), .IN2(n709), .QN(n708) );
  INVX0 U747 ( .INP(n706), .ZN(n566) );
  INVX0 U748 ( .INP(n709), .ZN(n684) );
  OA21X1 U749 ( .IN1(n710), .IN2(n711), .IN3(n712), .Q(n709) );
  XNOR2X1 U750 ( .IN1(n713), .IN2(keyinput38), .Q(n712) );
  NAND2X0 U751 ( .IN1(n711), .IN2(n710), .QN(n713) );
  XOR2X1 U752 ( .IN1(keyinput28), .IN2(n714), .Q(n711) );
  OA21X1 U753 ( .IN1(n481), .IN2(n715), .IN3(n716), .Q(n714) );
  XOR2X1 U754 ( .IN1(keyinput15), .IN2(n717), .Q(n716) );
  NOR2X0 U755 ( .IN1(n718), .IN2(n715), .QN(n717) );
  INVX0 U756 ( .INP(G6), .ZN(n718) );
  XNOR2X1 U757 ( .IN1(n719), .IN2(keyinput6), .Q(n715) );
  NAND2X0 U758 ( .IN1(G6), .IN2(G5), .QN(n719) );
  INVX0 U759 ( .INP(G5), .ZN(n481) );
  XNOR3X1 U760 ( .IN1(keyinput29), .IN2(G8), .IN3(n475), .Q(n710) );
  INVX0 U761 ( .INP(G7), .ZN(n475) );
  NAND2X0 U762 ( .IN1(n720), .IN2(n721), .QN(n706) );
  NAND3X0 U763 ( .IN1(n722), .IN2(n723), .IN3(n724), .QN(n721) );
  XOR2X1 U764 ( .IN1(keyinput37), .IN2(n725), .Q(n720) );
  AOI21X1 U765 ( .IN1(n723), .IN2(n722), .IN3(n724), .QN(n725) );
  XOR2X1 U766 ( .IN1(n726), .IN2(keyinput27), .Q(n724) );
  NAND2X0 U767 ( .IN1(n727), .IN2(n728), .QN(n726) );
  XOR2X1 U768 ( .IN1(n729), .IN2(keyinput13), .Q(n728) );
  OR2X1 U769 ( .IN1(n556), .IN2(G4), .Q(n729) );
  XOR2X1 U770 ( .IN1(n730), .IN2(keyinput14), .Q(n727) );
  NAND2X0 U771 ( .IN1(G4), .IN2(n556), .QN(n730) );
  INVX0 U772 ( .INP(G3), .ZN(n556) );
  XNOR2X1 U773 ( .IN1(n731), .IN2(keyinput5), .Q(n722) );
  NAND2X0 U774 ( .IN1(G2), .IN2(G1), .QN(n731) );
  OR2X1 U775 ( .IN1(G2), .IN2(G1), .Q(n723) );
  XOR3X1 U776 ( .IN1(keyinput45), .IN2(keyinput3), .IN3(n732), .Q(n693) );
  XNOR2X1 U777 ( .IN1(keyinput60), .IN2(keyinput52), .Q(n732) );
  XOR2X1 U778 ( .IN1(keyinput71), .IN2(n496), .Q(n560) );
  INVX0 U779 ( .INP(n413), .ZN(n496) );
  AO21X1 U780 ( .IN1(n733), .IN2(n734), .IN3(n735), .Q(n413) );
  XOR2X1 U781 ( .IN1(keyinput66), .IN2(n736), .Q(n735) );
  AND2X1 U782 ( .IN1(n733), .IN2(n737), .Q(n736) );
  XNOR2X1 U783 ( .IN1(n738), .IN2(keyinput61), .Q(n733) );
  NAND2X0 U784 ( .IN1(n737), .IN2(n734), .QN(n738) );
  AO21X1 U785 ( .IN1(n739), .IN2(n740), .IN3(n741), .Q(n734) );
  XOR2X1 U786 ( .IN1(keyinput42), .IN2(n742), .Q(n741) );
  NOR2X0 U787 ( .IN1(n743), .IN2(n744), .QN(n742) );
  INVX0 U788 ( .INP(n739), .ZN(n744) );
  XOR2X1 U789 ( .IN1(n640), .IN2(G22), .Q(n743) );
  INVX0 U790 ( .INP(G18), .ZN(n640) );
  XOR2X1 U791 ( .IN1(n745), .IN2(keyinput36), .Q(n739) );
  NAND2X0 U792 ( .IN1(n746), .IN2(n740), .QN(n745) );
  AO21X1 U793 ( .IN1(G26), .IN2(n409), .IN3(n747), .Q(n740) );
  XOR2X1 U794 ( .IN1(n748), .IN2(keyinput26), .Q(n747) );
  NAND2X0 U795 ( .IN1(G30), .IN2(n421), .QN(n748) );
  INVX0 U796 ( .INP(G26), .ZN(n421) );
  INVX0 U797 ( .INP(G30), .ZN(n409) );
  XOR2X1 U798 ( .IN1(G22), .IN2(G18), .Q(n746) );
  XOR3X1 U799 ( .IN1(n567), .IN2(n749), .IN3(n687), .Q(n737) );
  AO22X1 U800 ( .IN1(n750), .IN2(n751), .IN3(keyinput39), .IN4(n752), .Q(n687)
         );
  NAND2X0 U801 ( .IN1(n753), .IN2(n751), .QN(n752) );
  NAND2X0 U802 ( .IN1(n754), .IN2(n753), .QN(n751) );
  AO21X1 U803 ( .IN1(n753), .IN2(n755), .IN3(n754), .Q(n750) );
  XOR2X1 U804 ( .IN1(G14), .IN2(G13), .Q(n754) );
  INVX0 U805 ( .INP(keyinput39), .ZN(n755) );
  AO21X1 U806 ( .IN1(G15), .IN2(n673), .IN3(n756), .Q(n753) );
  XOR2X1 U807 ( .IN1(n757), .IN2(keyinput17), .Q(n756) );
  NAND2X0 U808 ( .IN1(G16), .IN2(n652), .QN(n757) );
  INVX0 U809 ( .INP(G15), .ZN(n652) );
  INVX0 U810 ( .INP(G16), .ZN(n673) );
  XNOR2X1 U811 ( .IN1(n758), .IN2(keyinput4), .Q(n749) );
  NAND2X0 U812 ( .IN1(G38), .IN2(G41), .QN(n758) );
  XOR3X1 U813 ( .IN1(keyinput44), .IN2(n468), .IN3(n759), .Q(n567) );
  XNOR2X1 U814 ( .IN1(G10), .IN2(n760), .Q(n759) );
  OA21X1 U815 ( .IN1(G11), .IN2(n672), .IN3(n761), .Q(n760) );
  XOR2X1 U816 ( .IN1(n762), .IN2(keyinput16), .Q(n761) );
  NAND2X0 U817 ( .IN1(G11), .IN2(n672), .QN(n762) );
  INVX0 U818 ( .INP(G12), .ZN(n672) );
  INVX0 U819 ( .INP(G9), .ZN(n468) );
endmodule

