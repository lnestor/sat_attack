
module c2670 ( N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, 
        N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, 
        N37, N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, 
        N57, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, 
        N75, N76, N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, 
        N91, N92, N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, 
        N106, N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119, 
        N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N135, 
        N136, N137, N138, N139, N140, N141, N142, N219, N224, N227, N230, N231, 
        N234, N237, N241, N246, N253, N256, N259, N262, N263, N266, N269, N272, 
        N275, N278, N281, N284, N287, N290, N294, N297, N301, N305, N309, N313, 
        N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, 
        N352, N355, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I, N149_I, 
        N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I, N157_I, N158_I, 
        N159_I, N160_I, N161_I, N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, 
        N168_I, N169_I, N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, 
        N177_I, N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I, 
        N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, 
        N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, 
        N204_I, N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I, 
        N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N398, N400, N401, N419, 
        N420, N456, N457, N458, N487, N488, N489, N490, N491, N492, N493, N494, 
        N792, N799, N805, N1026, N1028, N1029, N1269, N1277, N1448, N1726, 
        N1816, N1817, N1818, N1819, N1820, N1821, N1969, N1970, N1971, N2010, 
        N2012, N2014, N2016, N2018, N2020, N2022, N2387, N2388, N2389, N2390, 
        N2496, N2643, N2644, N2891, N2925, N2970, N2971, N3038, N3079, N3546, 
        N3671, N3803, N3804, N3809, N3851, N3875, N3881, N3882, N143_O, N144_O, 
        N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, N151_O, N152_O, N153_O, 
        N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, N160_O, N161_O, N162_O, 
        N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, 
        N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, 
        N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O, 
        N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O, N198_O, 
        N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O, N206_O, N207_O, 
        N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, N214_O, N215_O, N216_O, 
        N217_O, N218_O, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22,
         N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40,
         N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76,
         N77, N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N99, N100, N101, N102, N103, N104, N105, N106,
         N107, N108, N111, N112, N113, N114, N115, N116, N117, N118, N119,
         N120, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N135, N136, N137, N138, N139, N140, N141, N142, N219, N224, N227,
         N230, N231, N234, N237, N241, N246, N253, N256, N259, N262, N263,
         N266, N269, N272, N275, N278, N281, N284, N287, N290, N294, N297,
         N301, N305, N309, N313, N316, N319, N322, N325, N328, N331, N334,
         N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, N145_I,
         N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I,
         N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I,
         N162_I, N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I,
         N170_I, N171_I, N172_I, N173_I, N174_I, N175_I, N176_I, N177_I,
         N178_I, N179_I, N180_I, N181_I, N182_I, N183_I, N184_I, N185_I,
         N186_I, N187_I, N188_I, N189_I, N190_I, N191_I, N192_I, N193_I,
         N194_I, N195_I, N196_I, N197_I, N198_I, N199_I, N200_I, N201_I,
         N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, N208_I, N209_I,
         N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, N217_I,
         N218_I, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
         keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10,
         keyinput11, keyinput12, keyinput13, keyinput14, keyinput15,
         keyinput16, keyinput17, keyinput18, keyinput19, keyinput20,
         keyinput21, keyinput22, keyinput23, keyinput24, keyinput25,
         keyinput26, keyinput27, keyinput28, keyinput29, keyinput30,
         keyinput31, keyinput32, keyinput33, keyinput34, keyinput35,
         keyinput36, keyinput37, keyinput38, keyinput39, keyinput40,
         keyinput41, keyinput42, keyinput43, keyinput44, keyinput45,
         keyinput46, keyinput47, keyinput48, keyinput49, keyinput50,
         keyinput51, keyinput52, keyinput53, keyinput54, keyinput55,
         keyinput56, keyinput57, keyinput58, keyinput59, keyinput60,
         keyinput61, keyinput62, keyinput63, keyinput64, keyinput65,
         keyinput66, keyinput67, keyinput68, keyinput69, keyinput70,
         keyinput71, keyinput72, keyinput73, keyinput74, keyinput75,
         keyinput76, keyinput77, keyinput78, keyinput79, keyinput80,
         keyinput81, keyinput82, keyinput83, keyinput84, keyinput85,
         keyinput86, keyinput87, keyinput88, keyinput89, keyinput90,
         keyinput91, keyinput92, keyinput93, keyinput94, keyinput95,
         keyinput96, keyinput97, keyinput98, keyinput99, keyinput100,
         keyinput101, keyinput102, keyinput103, keyinput104, keyinput105,
         keyinput106, keyinput107, keyinput108, keyinput109, keyinput110,
         keyinput111, keyinput112, keyinput113, keyinput114, keyinput115,
         keyinput116, keyinput117, keyinput118, keyinput119, keyinput120,
         keyinput121, keyinput122, keyinput123, keyinput124, keyinput125,
         keyinput126, keyinput127;
  output N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489,
         N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029,
         N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821,
         N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022,
         N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970,
         N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875,
         N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O,
         N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O,
         N158_O, N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O,
         N166_O, N167_O, N168_O, N169_O, N170_O, N171_O, N172_O, N173_O,
         N174_O, N175_O, N176_O, N177_O, N178_O, N179_O, N180_O, N181_O,
         N182_O, N183_O, N184_O, N185_O, N186_O, N187_O, N188_O, N189_O,
         N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, N196_O, N197_O,
         N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, N205_O,
         N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O,
         N214_O, N215_O, N216_O, N217_O, N218_O;
  wire   N219, N253, N290, N143_I, N144_I, N145_I, N146_I, N147_I, N148_I,
         N149_I, N150_I, N151_I, N152_I, N153_I, N154_I, N155_I, N156_I,
         N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, N163_I, N164_I,
         N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, N172_I,
         N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I,
         N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I,
         N189_I, N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I,
         N197_I, N198_I, N199_I, N200_I, N201_I, N202_I, N203_I, N204_I,
         N205_I, N206_I, N207_I, N208_I, N209_I, N210_I, N211_I, N212_I,
         N213_I, N214_I, N215_I, N216_I, N217_I, N218_I, N2387, N2389, N2643,
         N3803, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994;
  assign N805 = N219;
  assign N401 = N219;
  assign N400 = N219;
  assign N398 = N219;
  assign N420 = N253;
  assign N419 = N253;
  assign N458 = N290;
  assign N457 = N290;
  assign N456 = N290;
  assign N143_O = N143_I;
  assign N144_O = N144_I;
  assign N145_O = N145_I;
  assign N146_O = N146_I;
  assign N147_O = N147_I;
  assign N148_O = N148_I;
  assign N149_O = N149_I;
  assign N150_O = N150_I;
  assign N151_O = N151_I;
  assign N152_O = N152_I;
  assign N153_O = N153_I;
  assign N154_O = N154_I;
  assign N155_O = N155_I;
  assign N156_O = N156_I;
  assign N157_O = N157_I;
  assign N158_O = N158_I;
  assign N159_O = N159_I;
  assign N160_O = N160_I;
  assign N161_O = N161_I;
  assign N162_O = N162_I;
  assign N163_O = N163_I;
  assign N164_O = N164_I;
  assign N165_O = N165_I;
  assign N166_O = N166_I;
  assign N167_O = N167_I;
  assign N168_O = N168_I;
  assign N169_O = N169_I;
  assign N170_O = N170_I;
  assign N171_O = N171_I;
  assign N172_O = N172_I;
  assign N173_O = N173_I;
  assign N174_O = N174_I;
  assign N175_O = N175_I;
  assign N176_O = N176_I;
  assign N177_O = N177_I;
  assign N178_O = N178_I;
  assign N179_O = N179_I;
  assign N180_O = N180_I;
  assign N181_O = N181_I;
  assign N182_O = N182_I;
  assign N183_O = N183_I;
  assign N184_O = N184_I;
  assign N185_O = N185_I;
  assign N186_O = N186_I;
  assign N187_O = N187_I;
  assign N188_O = N188_I;
  assign N189_O = N189_I;
  assign N190_O = N190_I;
  assign N191_O = N191_I;
  assign N192_O = N192_I;
  assign N193_O = N193_I;
  assign N194_O = N194_I;
  assign N195_O = N195_I;
  assign N196_O = N196_I;
  assign N197_O = N197_I;
  assign N198_O = N198_I;
  assign N199_O = N199_I;
  assign N200_O = N200_I;
  assign N201_O = N201_I;
  assign N202_O = N202_I;
  assign N203_O = N203_I;
  assign N204_O = N204_I;
  assign N205_O = N205_I;
  assign N206_O = N206_I;
  assign N207_O = N207_I;
  assign N208_O = N208_I;
  assign N209_O = N209_I;
  assign N210_O = N210_I;
  assign N211_O = N211_I;
  assign N212_O = N212_I;
  assign N213_O = N213_I;
  assign N214_O = N214_I;
  assign N215_O = N215_I;
  assign N216_O = N216_I;
  assign N217_O = N217_I;
  assign N218_O = N218_I;
  assign N2388 = N2387;
  assign N2390 = N2389;
  assign N2644 = N2643;
  assign N3804 = N3803;

  XOR2X1 U540 ( .IN1(n520), .IN2(keyinput3), .Q(N799) );
  NAND3X0 U541 ( .IN1(N2), .IN2(N15), .IN3(N237), .QN(n520) );
  XNOR2X1 U542 ( .IN1(n521), .IN2(keyinput9), .Q(N792) );
  NAND4X0 U543 ( .IN1(N309), .IN2(N305), .IN3(N301), .IN4(N297), .QN(n521) );
  INVX0 U544 ( .INP(N108), .ZN(N494) );
  XNOR2X1 U545 ( .IN1(N57), .IN2(keyinput2), .Q(N493) );
  INVX0 U546 ( .INP(N120), .ZN(N492) );
  INVX0 U547 ( .INP(N69), .ZN(N491) );
  INVX0 U548 ( .INP(N96), .ZN(N490) );
  INVX0 U549 ( .INP(N82), .ZN(N489) );
  INVX0 U550 ( .INP(N132), .ZN(N488) );
  XOR2X1 U551 ( .IN1(keyinput1), .IN2(N44), .Q(N487) );
  INVX0 U552 ( .INP(N3882), .ZN(N3881) );
  NAND4X0 U553 ( .IN1(n522), .IN2(n523), .IN3(N1726), .IN4(n524), .QN(N3882)
         );
  NOR4X0 U554 ( .IN1(N3875), .IN2(N3809), .IN3(N3671), .IN4(N2925), .QN(n524)
         );
  INVX0 U555 ( .INP(N2971), .ZN(n523) );
  INVX0 U556 ( .INP(N2970), .ZN(n522) );
  AND2X1 U557 ( .IN1(keyinput127), .IN2(n525), .Q(N3875) );
  XOR2X1 U558 ( .IN1(keyinput126), .IN2(n526), .Q(n525) );
  OA21X1 U559 ( .IN1(N3851), .IN2(n527), .IN3(n528), .Q(n526) );
  XOR2X1 U560 ( .IN1(n529), .IN2(keyinput125), .Q(n528) );
  NAND2X0 U561 ( .IN1(n527), .IN2(N3851), .QN(n529) );
  XNOR2X1 U562 ( .IN1(keyinput124), .IN2(n530), .Q(n527) );
  OA222X1 U563 ( .IN1(n531), .IN2(n532), .IN3(n533), .IN4(n534), .IN5(n535), 
        .IN6(n536), .Q(n530) );
  INVX0 U564 ( .INP(n537), .ZN(n536) );
  OA21X1 U565 ( .IN1(n538), .IN2(n539), .IN3(n540), .Q(n535) );
  NAND3X0 U566 ( .IN1(n541), .IN2(n542), .IN3(n543), .QN(n540) );
  AO222X1 U567 ( .IN1(n544), .IN2(n545), .IN3(n546), .IN4(n547), .IN5(n548), 
        .IN6(n549), .Q(n541) );
  INVX0 U568 ( .INP(n550), .ZN(n548) );
  AND2X1 U569 ( .IN1(n533), .IN2(n551), .Q(n546) );
  INVX0 U570 ( .INP(n552), .ZN(n539) );
  NAND2X0 U571 ( .IN1(n553), .IN2(n547), .QN(n534) );
  OAI22X1 U572 ( .IN1(n554), .IN2(n555), .IN3(n556), .IN4(n557), .QN(n547) );
  OA21X1 U573 ( .IN1(keyinput109), .IN2(n554), .IN3(n555), .Q(n556) );
  XOR2X1 U574 ( .IN1(n558), .IN2(keyinput88), .Q(n555) );
  NAND2X0 U575 ( .IN1(n559), .IN2(N2020), .QN(n558) );
  OA21X1 U576 ( .IN1(n560), .IN2(n561), .IN3(n562), .Q(n554) );
  XOR2X1 U577 ( .IN1(n563), .IN2(keyinput103), .Q(n562) );
  NAND2X0 U578 ( .IN1(n564), .IN2(n565), .QN(n563) );
  OA21X1 U579 ( .IN1(n564), .IN2(n566), .IN3(n567), .Q(n561) );
  XOR2X1 U580 ( .IN1(n568), .IN2(keyinput112), .Q(n567) );
  NAND2X0 U581 ( .IN1(n566), .IN2(n564), .QN(n568) );
  INVX0 U582 ( .INP(n565), .ZN(n566) );
  NAND2X0 U583 ( .IN1(n559), .IN2(N2018), .QN(n565) );
  NOR2X0 U584 ( .IN1(n569), .IN2(n570), .QN(n559) );
  OA22X1 U585 ( .IN1(n571), .IN2(n572), .IN3(n573), .IN4(n574), .Q(n560) );
  AND2X1 U586 ( .IN1(n574), .IN2(n573), .Q(n572) );
  AOI21X1 U587 ( .IN1(n570), .IN2(n575), .IN3(n576), .QN(n573) );
  AOI21X1 U588 ( .IN1(n577), .IN2(n578), .IN3(n579), .QN(n574) );
  OA22X1 U589 ( .IN1(n577), .IN2(n578), .IN3(n580), .IN4(n581), .Q(n579) );
  NOR2X0 U590 ( .IN1(n582), .IN2(n583), .QN(n580) );
  OA22X1 U591 ( .IN1(n584), .IN2(n585), .IN3(N2010), .IN4(n586), .Q(n582) );
  INVX0 U592 ( .INP(n587), .ZN(n586) );
  OA21X1 U593 ( .IN1(n588), .IN2(n589), .IN3(n590), .Q(n585) );
  NAND3X0 U594 ( .IN1(n591), .IN2(n592), .IN3(n593), .QN(n590) );
  XNOR2X1 U595 ( .IN1(n594), .IN2(keyinput102), .Q(n593) );
  AO21X1 U596 ( .IN1(keyinput68), .IN2(n595), .IN3(n596), .Q(n592) );
  INVX0 U597 ( .INP(n595), .ZN(n588) );
  AO21X1 U598 ( .IN1(n597), .IN2(n598), .IN3(n599), .Q(n595) );
  XOR2X1 U599 ( .IN1(n600), .IN2(keyinput90), .Q(n599) );
  NAND2X0 U600 ( .IN1(n601), .IN2(n575), .QN(n600) );
  NOR2X0 U601 ( .IN1(n602), .IN2(n587), .QN(n584) );
  MUX21X1 U602 ( .IN1(n603), .IN2(n604), .S(n575), .Q(n587) );
  AO21X1 U603 ( .IN1(n605), .IN2(n606), .IN3(n607), .Q(n578) );
  NAND3X0 U604 ( .IN1(n608), .IN2(N2014), .IN3(N8), .QN(n577) );
  NAND2X0 U605 ( .IN1(n570), .IN2(n575), .QN(n608) );
  XNOR2X1 U606 ( .IN1(n597), .IN2(keyinput78), .Q(n570) );
  NAND4X0 U607 ( .IN1(n543), .IN2(n537), .IN3(n551), .IN4(n542), .QN(n553) );
  NAND3X0 U608 ( .IN1(n609), .IN2(n610), .IN3(n538), .QN(n542) );
  NAND2X0 U609 ( .IN1(keyinput108), .IN2(n552), .QN(n610) );
  OR3X1 U610 ( .IN1(n545), .IN2(n544), .IN3(n611), .Q(n551) );
  NAND2X0 U611 ( .IN1(n531), .IN2(n612), .QN(n537) );
  XNOR2X1 U612 ( .IN1(keyinput111), .IN2(n532), .Q(n612) );
  NAND2X0 U613 ( .IN1(n613), .IN2(n550), .QN(n543) );
  NAND2X0 U614 ( .IN1(n609), .IN2(n614), .QN(n550) );
  XNOR2X1 U615 ( .IN1(keyinput92), .IN2(n615), .Q(n614) );
  INVX0 U616 ( .INP(n549), .ZN(n613) );
  NAND2X0 U617 ( .IN1(n616), .IN2(n609), .QN(n549) );
  XOR2X1 U618 ( .IN1(n617), .IN2(keyinput73), .Q(n616) );
  INVX0 U619 ( .INP(keyinput116), .ZN(n533) );
  INVX0 U620 ( .INP(n618), .ZN(n532) );
  AND2X1 U621 ( .IN1(n619), .IN2(n609), .Q(n531) );
  XNOR2X1 U622 ( .IN1(n620), .IN2(keyinput74), .Q(n619) );
  NAND2X0 U623 ( .IN1(n621), .IN2(n622), .QN(N3851) );
  NAND4X0 U624 ( .IN1(n623), .IN2(n624), .IN3(n625), .IN4(n626), .QN(n622) );
  OA21X1 U625 ( .IN1(n627), .IN2(n628), .IN3(n629), .Q(n625) );
  XOR2X1 U626 ( .IN1(n630), .IN2(keyinput123), .Q(n624) );
  NAND2X0 U627 ( .IN1(n631), .IN2(n632), .QN(n630) );
  XNOR2X1 U628 ( .IN1(keyinput121), .IN2(n633), .Q(n632) );
  OA221X1 U629 ( .IN1(n634), .IN2(n635), .IN3(n636), .IN4(keyinput118), .IN5(
        n637), .Q(n633) );
  INVX0 U630 ( .INP(n638), .ZN(n637) );
  NOR4X0 U631 ( .IN1(n639), .IN2(n571), .IN3(n635), .IN4(n640), .QN(n636) );
  OA21X1 U632 ( .IN1(n641), .IN2(n640), .IN3(n642), .Q(n634) );
  OA22X1 U633 ( .IN1(n643), .IN2(n644), .IN3(n645), .IN4(n646), .Q(n641) );
  OA21X1 U634 ( .IN1(n647), .IN2(n648), .IN3(n649), .Q(n645) );
  INVX0 U635 ( .INP(n650), .ZN(n649) );
  NAND2X0 U636 ( .IN1(n651), .IN2(n576), .QN(n644) );
  INVX0 U637 ( .INP(n639), .ZN(n576) );
  INVX0 U638 ( .INP(keyinput118), .ZN(n643) );
  XNOR2X1 U639 ( .IN1(keyinput122), .IN2(n652), .Q(n631) );
  NOR2X0 U640 ( .IN1(n653), .IN2(n654), .QN(n652) );
  XOR2X1 U641 ( .IN1(n655), .IN2(keyinput120), .Q(n654) );
  OR4X1 U642 ( .IN1(n640), .IN2(n635), .IN3(n647), .IN4(n656), .Q(n655) );
  OR2X1 U643 ( .IN1(n583), .IN2(n646), .Q(n656) );
  XNOR2X1 U644 ( .IN1(n657), .IN2(n639), .Q(n646) );
  NOR2X0 U645 ( .IN1(n569), .IN2(N1819), .QN(n639) );
  NAND2X0 U646 ( .IN1(keyinput113), .IN2(n651), .QN(n657) );
  INVX0 U647 ( .INP(n571), .ZN(n651) );
  OA22X1 U648 ( .IN1(n658), .IN2(N272), .IN3(n659), .IN4(n575), .Q(n571) );
  OR2X1 U649 ( .IN1(N309), .IN2(n569), .Q(n659) );
  AO21X1 U650 ( .IN1(n660), .IN2(n661), .IN3(n581), .Q(n583) );
  INVX0 U651 ( .INP(n648), .ZN(n581) );
  NAND2X0 U652 ( .IN1(n662), .IN2(n663), .QN(n648) );
  MUX21X1 U653 ( .IN1(n664), .IN2(n665), .S(n575), .Q(n662) );
  INVX0 U654 ( .INP(n663), .ZN(n661) );
  MUX21X1 U655 ( .IN1(N301), .IN2(N266), .S(n575), .Q(n660) );
  AO21X1 U656 ( .IN1(n666), .IN2(n667), .IN3(n650), .Q(n647) );
  NOR2X0 U657 ( .IN1(n667), .IN2(n666), .QN(n650) );
  AO22X1 U658 ( .IN1(n605), .IN2(N2014), .IN3(n668), .IN4(N8), .Q(n667) );
  XNOR2X1 U659 ( .IN1(N1820), .IN2(keyinput76), .Q(n668) );
  XOR2X1 U660 ( .IN1(keyinput110), .IN2(n669), .Q(n666) );
  NOR2X0 U661 ( .IN1(n607), .IN2(n670), .QN(n669) );
  MUX21X1 U662 ( .IN1(n671), .IN2(n672), .S(keyinput93), .Q(n670) );
  OA21X1 U663 ( .IN1(n597), .IN2(N269), .IN3(N8), .Q(n672) );
  NOR2X0 U664 ( .IN1(N269), .IN2(n658), .QN(n671) );
  AND3X1 U665 ( .IN1(N8), .IN2(n673), .IN3(n597), .Q(n607) );
  AO21X1 U666 ( .IN1(n674), .IN2(n557), .IN3(n638), .Q(n635) );
  NOR2X0 U667 ( .IN1(n557), .IN2(n674), .QN(n638) );
  NAND2X0 U668 ( .IN1(n605), .IN2(n675), .QN(n557) );
  NOR2X0 U669 ( .IN1(n658), .IN2(n676), .QN(n674) );
  NAND2X0 U670 ( .IN1(n642), .IN2(n677), .QN(n640) );
  OR3X1 U671 ( .IN1(n678), .IN2(n564), .IN3(n658), .Q(n677) );
  NAND2X0 U672 ( .IN1(n564), .IN2(n678), .QN(n642) );
  NOR2X0 U673 ( .IN1(n658), .IN2(N275), .QN(n564) );
  INVX0 U674 ( .INP(n605), .ZN(n658) );
  NOR2X0 U675 ( .IN1(n569), .IN2(n597), .QN(n605) );
  INVX0 U676 ( .INP(N8), .ZN(n569) );
  OA22X1 U677 ( .IN1(N2010), .IN2(n679), .IN3(n680), .IN4(n681), .Q(n653) );
  AND2X1 U678 ( .IN1(n681), .IN2(n680), .Q(n679) );
  AND2X1 U679 ( .IN1(n682), .IN2(n683), .Q(n680) );
  XOR2X1 U680 ( .IN1(n684), .IN2(keyinput101), .Q(n683) );
  NAND2X0 U681 ( .IN1(n597), .IN2(n603), .QN(n684) );
  XOR2X1 U682 ( .IN1(n685), .IN2(keyinput91), .Q(n682) );
  NAND2X0 U683 ( .IN1(n604), .IN2(n575), .QN(n685) );
  AO21X1 U684 ( .IN1(n686), .IN2(n589), .IN3(n687), .Q(n681) );
  OA22X1 U685 ( .IN1(n686), .IN2(n589), .IN3(n594), .IN4(n688), .Q(n687) );
  MUX21X1 U686 ( .IN1(N287), .IN2(N256), .S(n575), .Q(n594) );
  MUX21X1 U687 ( .IN1(N259), .IN2(N294), .S(n597), .Q(n686) );
  INVX0 U688 ( .INP(n575), .ZN(n597) );
  NAND4X0 U689 ( .IN1(n689), .IN2(N40), .IN3(N1816), .IN4(n690), .QN(n575) );
  XOR2X1 U690 ( .IN1(n691), .IN2(n544), .Q(n623) );
  XNOR2X1 U691 ( .IN1(n692), .IN2(keyinput119), .Q(n621) );
  NAND3X0 U692 ( .IN1(n693), .IN2(n694), .IN3(n695), .QN(n692) );
  XNOR2X1 U693 ( .IN1(n696), .IN2(keyinput117), .Q(n695) );
  NAND3X0 U694 ( .IN1(n697), .IN2(n698), .IN3(n626), .QN(n696) );
  NAND3X0 U695 ( .IN1(n629), .IN2(n699), .IN3(n626), .QN(n693) );
  OA21X1 U696 ( .IN1(n700), .IN2(n618), .IN3(n694), .Q(n626) );
  NAND2X0 U697 ( .IN1(n618), .IN2(n700), .QN(n694) );
  NOR2X0 U698 ( .IN1(n611), .IN2(N294), .QN(n618) );
  NAND2X0 U699 ( .IN1(n701), .IN2(n609), .QN(n700) );
  XOR2X1 U700 ( .IN1(n702), .IN2(keyinput77), .Q(n701) );
  OR2X1 U701 ( .IN1(keyinput69), .IN2(n620), .Q(n702) );
  NAND2X0 U702 ( .IN1(n703), .IN2(n704), .QN(n699) );
  NAND3X0 U703 ( .IN1(n705), .IN2(n691), .IN3(n544), .QN(n704) );
  NOR2X0 U704 ( .IN1(n611), .IN2(N281), .QN(n544) );
  NAND2X0 U705 ( .IN1(n706), .IN2(N2022), .QN(n691) );
  OR2X1 U706 ( .IN1(n628), .IN2(n627), .Q(n705) );
  NOR2X0 U707 ( .IN1(n707), .IN2(n708), .QN(n627) );
  XOR2X1 U708 ( .IN1(n709), .IN2(keyinput114), .Q(n628) );
  NAND2X0 U709 ( .IN1(n707), .IN2(n708), .QN(n709) );
  XOR2X1 U710 ( .IN1(keyinput104), .IN2(n710), .Q(n703) );
  NOR2X0 U711 ( .IN1(n711), .IN2(n708), .QN(n710) );
  NAND2X0 U712 ( .IN1(n712), .IN2(n609), .QN(n708) );
  INVX0 U713 ( .INP(n611), .ZN(n609) );
  XNOR2X1 U714 ( .IN1(N284), .IN2(keyinput94), .Q(n712) );
  INVX0 U715 ( .INP(n707), .ZN(n711) );
  NAND2X0 U716 ( .IN1(n706), .IN2(n617), .QN(n707) );
  XOR2X1 U717 ( .IN1(n697), .IN2(n698), .Q(n629) );
  NAND2X0 U718 ( .IN1(n538), .IN2(n706), .QN(n698) );
  NOR2X0 U719 ( .IN1(n611), .IN2(keyinput69), .QN(n706) );
  XNOR2X1 U720 ( .IN1(n713), .IN2(keyinput98), .Q(n697) );
  MUX21X1 U721 ( .IN1(n552), .IN2(n714), .S(keyinput95), .Q(n713) );
  NOR2X0 U722 ( .IN1(n611), .IN2(n715), .QN(n714) );
  NOR2X0 U723 ( .IN1(n611), .IN2(N287), .QN(n552) );
  NAND3X0 U724 ( .IN1(N1816), .IN2(n716), .IN3(N40), .QN(n611) );
  NAND2X0 U725 ( .IN1(n689), .IN2(n690), .QN(n716) );
  XNOR2X1 U726 ( .IN1(N262), .IN2(keyinput0), .Q(n689) );
  AND2X1 U727 ( .IN1(n717), .IN2(n718), .Q(N3809) );
  XOR3X1 U728 ( .IN1(n719), .IN2(n720), .IN3(n721), .Q(n717) );
  NAND3X0 U729 ( .IN1(n722), .IN2(n723), .IN3(n724), .QN(n721) );
  XOR2X1 U730 ( .IN1(n725), .IN2(keyinput106), .Q(n724) );
  NAND2X0 U731 ( .IN1(n726), .IN2(n727), .QN(n725) );
  XOR2X1 U732 ( .IN1(n728), .IN2(n729), .Q(n727) );
  OR3X1 U733 ( .IN1(n728), .IN2(n726), .IN3(n729), .Q(n723) );
  INVX0 U734 ( .INP(n730), .ZN(n726) );
  XNOR2X1 U735 ( .IN1(n731), .IN2(keyinput100), .Q(n722) );
  NAND3X0 U736 ( .IN1(n729), .IN2(n730), .IN3(n728), .QN(n731) );
  XOR2X1 U737 ( .IN1(n663), .IN2(N1820), .Q(n728) );
  XOR2X1 U738 ( .IN1(N1821), .IN2(keyinput56), .Q(n663) );
  XNOR2X1 U739 ( .IN1(n602), .IN2(n589), .Q(n730) );
  XNOR2X1 U740 ( .IN1(n732), .IN2(N2016), .Q(n720) );
  NOR2X0 U741 ( .IN1(keyinput96), .IN2(n733), .QN(n732) );
  XNOR2X1 U742 ( .IN1(n545), .IN2(n734), .Q(n733) );
  MUX21X1 U743 ( .IN1(n735), .IN2(n736), .S(N246), .Q(N3803) );
  XOR2X1 U744 ( .IN1(n737), .IN2(n738), .Q(n736) );
  XOR3X1 U745 ( .IN1(n719), .IN2(n739), .IN3(n740), .Q(n738) );
  NAND2X0 U746 ( .IN1(n741), .IN2(keyinput107), .QN(n740) );
  MUX21X1 U747 ( .IN1(n742), .IN2(n743), .S(n729), .Q(n741) );
  XNOR2X1 U748 ( .IN1(n591), .IN2(n735), .Q(n729) );
  XNOR2X1 U749 ( .IN1(n744), .IN2(n745), .Q(n743) );
  NAND2X0 U750 ( .IN1(keyinput99), .IN2(n746), .QN(n744) );
  XOR2X1 U751 ( .IN1(n747), .IN2(n745), .Q(n742) );
  AO21X1 U752 ( .IN1(n596), .IN2(N2010), .IN3(n748), .Q(n745) );
  XOR2X1 U753 ( .IN1(keyinput75), .IN2(n749), .Q(n748) );
  NOR2X0 U754 ( .IN1(N2010), .IN2(n596), .QN(n749) );
  NAND2X0 U755 ( .IN1(keyinput83), .IN2(n734), .QN(n739) );
  XNOR2X1 U756 ( .IN1(N2020), .IN2(keyinput58), .Q(n734) );
  XNOR2X1 U757 ( .IN1(n678), .IN2(keyinput57), .Q(n719) );
  XNOR3X1 U758 ( .IN1(keyinput115), .IN2(n750), .IN3(n545), .Q(n737) );
  INVX0 U759 ( .INP(N2022), .ZN(n545) );
  NOR2X0 U760 ( .IN1(keyinput82), .IN2(N2016), .QN(n750) );
  AND2X1 U761 ( .IN1(n751), .IN2(n718), .Q(N3671) );
  INVX0 U762 ( .INP(N37), .ZN(n718) );
  XOR3X1 U763 ( .IN1(n752), .IN2(n753), .IN3(n754), .Q(n751) );
  XNOR3X1 U764 ( .IN1(n755), .IN2(n756), .IN3(n757), .Q(n754) );
  AO221X1 U765 ( .IN1(N106), .IN2(n758), .IN3(N118), .IN4(n759), .IN5(n760), 
        .Q(n756) );
  AO21X1 U766 ( .IN1(N130), .IN2(n761), .IN3(n762), .Q(n760) );
  XOR2X1 U767 ( .IN1(n763), .IN2(keyinput35), .Q(n762) );
  NAND2X0 U768 ( .IN1(N142), .IN2(n764), .QN(n763) );
  NOR2X0 U769 ( .IN1(keyinput81), .IN2(n765), .QN(n755) );
  XNOR2X1 U770 ( .IN1(n766), .IN2(n767), .Q(n765) );
  OA21X1 U771 ( .IN1(n768), .IN2(n690), .IN3(n769), .Q(n767) );
  XOR2X1 U772 ( .IN1(n770), .IN2(keyinput63), .Q(n769) );
  NAND2X0 U773 ( .IN1(n768), .IN2(n690), .QN(n770) );
  OA21X1 U774 ( .IN1(n771), .IN2(n772), .IN3(n773), .Q(n766) );
  XOR2X1 U775 ( .IN1(keyinput62), .IN2(n774), .Q(n773) );
  NOR2X0 U776 ( .IN1(n620), .IN2(n538), .QN(n774) );
  XOR2X1 U777 ( .IN1(n617), .IN2(n775), .Q(n753) );
  XOR2X1 U778 ( .IN1(keyinput87), .IN2(n776), .Q(n752) );
  OA21X1 U779 ( .IN1(N1817), .IN2(n777), .IN3(n778), .Q(n776) );
  XOR2X1 U780 ( .IN1(keyinput66), .IN2(n779), .Q(n778) );
  NOR2X0 U781 ( .IN1(N1816), .IN2(n780), .QN(n779) );
  MUX21X1 U782 ( .IN1(n781), .IN2(n782), .S(n783), .Q(N2971) );
  MUX21X1 U783 ( .IN1(n784), .IN2(n785), .S(n786), .Q(n783) );
  XNOR2X1 U784 ( .IN1(N352), .IN2(n604), .Q(n786) );
  XOR2X1 U785 ( .IN1(n787), .IN2(n788), .Q(n785) );
  NOR2X0 U786 ( .IN1(keyinput53), .IN2(n789), .QN(n787) );
  XOR2X1 U787 ( .IN1(n789), .IN2(n788), .Q(n784) );
  XNOR2X1 U788 ( .IN1(n790), .IN2(N272), .Q(n788) );
  AO21X1 U789 ( .IN1(N266), .IN2(n606), .IN3(n791), .Q(n789) );
  XOR2X1 U790 ( .IN1(n792), .IN2(keyinput24), .Q(n791) );
  NAND2X0 U791 ( .IN1(N269), .IN2(n793), .QN(n792) );
  XNOR2X1 U792 ( .IN1(keyinput16), .IN2(n665), .Q(n793) );
  NAND2X0 U793 ( .IN1(n794), .IN2(n795), .QN(n782) );
  AND2X1 U794 ( .IN1(n795), .IN2(n794), .Q(n781) );
  XNOR2X1 U795 ( .IN1(n796), .IN2(keyinput52), .Q(n794) );
  OR2X1 U796 ( .IN1(n797), .IN2(n798), .Q(n796) );
  NAND2X0 U797 ( .IN1(n799), .IN2(n797), .QN(n795) );
  AO21X1 U798 ( .IN1(N281), .IN2(n675), .IN3(n800), .Q(n797) );
  XOR2X1 U799 ( .IN1(keyinput28), .IN2(n801), .Q(n800) );
  NOR2X0 U800 ( .IN1(N281), .IN2(n675), .QN(n801) );
  XOR2X1 U801 ( .IN1(keyinput46), .IN2(n798), .Q(n799) );
  XOR3X1 U802 ( .IN1(keyinput38), .IN2(n715), .IN3(n615), .Q(n798) );
  NAND2X0 U803 ( .IN1(n802), .IN2(n803), .QN(N3546) );
  AO21X1 U804 ( .IN1(n804), .IN2(keyinput47), .IN3(N241), .Q(n803) );
  XOR3X1 U805 ( .IN1(keyinput105), .IN2(n805), .IN3(n735), .Q(n804) );
  NOR2X0 U806 ( .IN1(keyinput67), .IN2(n806), .QN(n805) );
  XOR2X1 U807 ( .IN1(keyinput97), .IN2(n807), .Q(n806) );
  OA21X1 U808 ( .IN1(n746), .IN2(n808), .IN3(n809), .Q(n807) );
  XOR2X1 U809 ( .IN1(n810), .IN2(keyinput89), .Q(n809) );
  NAND2X0 U810 ( .IN1(n746), .IN2(n591), .QN(n810) );
  XNOR2X1 U811 ( .IN1(n596), .IN2(n591), .Q(n808) );
  MUX21X1 U812 ( .IN1(keyinput47), .IN2(n811), .S(n735), .Q(n802) );
  AO221X1 U813 ( .IN1(N80), .IN2(n812), .IN3(N67), .IN4(n813), .IN5(n814), .Q(
        n735) );
  AO22X1 U814 ( .IN1(N55), .IN2(n815), .IN3(N93), .IN4(n816), .Q(n814) );
  NAND2X0 U815 ( .IN1(keyinput47), .IN2(N241), .QN(n811) );
  INVX0 U816 ( .INP(N3038), .ZN(N3079) );
  NOR4X0 U817 ( .IN1(n817), .IN2(n818), .IN3(n819), .IN4(n820), .QN(N3038) );
  NAND4X0 U818 ( .IN1(n821), .IN2(n822), .IN3(n823), .IN4(n824), .QN(n820) );
  AND3X1 U819 ( .IN1(n825), .IN2(n826), .IN3(n827), .Q(n824) );
  XOR3X1 U820 ( .IN1(keyinput55), .IN2(n828), .IN3(n829), .Q(n827) );
  NAND2X0 U821 ( .IN1(keyinput65), .IN2(n715), .QN(n829) );
  INVX0 U822 ( .INP(N287), .ZN(n715) );
  MUX21X1 U823 ( .IN1(N32), .IN2(n538), .S(N29), .Q(n828) );
  INVX0 U824 ( .INP(n771), .ZN(n538) );
  XNOR2X1 U825 ( .IN1(n830), .IN2(keyinput42), .Q(n771) );
  AO221X1 U826 ( .IN1(N117), .IN2(n759), .IN3(N129), .IN4(n761), .IN5(n831), 
        .Q(n830) );
  AO22X1 U827 ( .IN1(N105), .IN2(n758), .IN3(N141), .IN4(n764), .Q(n831) );
  XNOR3X1 U828 ( .IN1(keyinput80), .IN2(n604), .IN3(n832), .Q(n826) );
  NOR2X0 U829 ( .IN1(n833), .IN2(keyinput34), .QN(n832) );
  OA21X1 U830 ( .IN1(n602), .IN2(n834), .IN3(n835), .Q(n833) );
  XOR2X1 U831 ( .IN1(n836), .IN2(keyinput37), .Q(n835) );
  NAND2X0 U832 ( .IN1(N20), .IN2(n834), .QN(n836) );
  INVX0 U833 ( .INP(N2010), .ZN(n602) );
  INVX0 U834 ( .INP(N263), .ZN(n604) );
  XNOR3X1 U835 ( .IN1(keyinput54), .IN2(n606), .IN3(n837), .Q(n825) );
  MUX21X1 U836 ( .IN1(N2014), .IN2(N21), .S(n834), .Q(n837) );
  INVX0 U837 ( .INP(N269), .ZN(n606) );
  XNOR2X1 U838 ( .IN1(n838), .IN2(n673), .Q(n823) );
  XOR2X1 U839 ( .IN1(N305), .IN2(keyinput8), .Q(n673) );
  AO22X1 U840 ( .IN1(N29), .IN2(n777), .IN3(N34), .IN4(n839), .Q(n838) );
  OR2X1 U841 ( .IN1(n775), .IN2(n840), .Q(n822) );
  XNOR2X1 U842 ( .IN1(n841), .IN2(keyinput85), .Q(n821) );
  NAND4X0 U843 ( .IN1(n842), .IN2(n843), .IN3(n844), .IN4(n845), .QN(n841) );
  OA221X1 U844 ( .IN1(n615), .IN2(n846), .IN3(N272), .IN4(n847), .IN5(n848), 
        .Q(n845) );
  NOR2X0 U845 ( .IN1(n849), .IN2(n850), .QN(n848) );
  XOR2X1 U846 ( .IN1(n851), .IN2(keyinput60), .Q(n850) );
  NAND2X0 U847 ( .IN1(N272), .IN2(n847), .QN(n851) );
  XNOR2X1 U848 ( .IN1(n852), .IN2(n853), .Q(n849) );
  NAND2X0 U849 ( .IN1(keyinput61), .IN2(n790), .QN(n853) );
  INVX0 U850 ( .INP(N275), .ZN(n790) );
  AO21X1 U851 ( .IN1(N23), .IN2(n834), .IN3(n854), .Q(n852) );
  XOR2X1 U852 ( .IN1(keyinput51), .IN2(n855), .Q(n854) );
  NOR2X0 U853 ( .IN1(n678), .IN2(n834), .QN(n855) );
  INVX0 U854 ( .INP(N2018), .ZN(n678) );
  AO21X1 U855 ( .IN1(N22), .IN2(n834), .IN3(n856), .Q(n847) );
  XOR2X1 U856 ( .IN1(n857), .IN2(keyinput50), .Q(n856) );
  NAND2X0 U857 ( .IN1(N16), .IN2(N2016), .QN(n857) );
  XNOR3X1 U858 ( .IN1(keyinput72), .IN2(n858), .IN3(N281), .Q(n844) );
  MUX21X1 U859 ( .IN1(N2022), .IN2(N24), .S(n834), .Q(n858) );
  XNOR2X1 U860 ( .IN1(keyinput79), .IN2(n859), .Q(n843) );
  OA21X1 U861 ( .IN1(n675), .IN2(n860), .IN3(n861), .Q(n859) );
  XOR2X1 U862 ( .IN1(n862), .IN2(keyinput70), .Q(n861) );
  NAND2X0 U863 ( .IN1(n860), .IN2(n675), .QN(n862) );
  MUX21X1 U864 ( .IN1(n676), .IN2(n863), .S(n834), .Q(n860) );
  INVX0 U865 ( .INP(N6), .ZN(n863) );
  INVX0 U866 ( .INP(N2020), .ZN(n676) );
  INVX0 U867 ( .INP(N278), .ZN(n675) );
  XOR2X1 U868 ( .IN1(n864), .IN2(keyinput71), .Q(n842) );
  NAND2X0 U869 ( .IN1(n846), .IN2(n615), .QN(n864) );
  INVX0 U870 ( .INP(N284), .ZN(n615) );
  INVX0 U871 ( .INP(n865), .ZN(n846) );
  MUX21X1 U872 ( .IN1(N25), .IN2(n617), .S(N29), .Q(n865) );
  AO221X1 U873 ( .IN1(N107), .IN2(n759), .IN3(N119), .IN4(n761), .IN5(n866), 
        .Q(n617) );
  AO22X1 U874 ( .IN1(N95), .IN2(n758), .IN3(N131), .IN4(n764), .Q(n866) );
  NAND3X0 U875 ( .IN1(n867), .IN2(n868), .IN3(n869), .QN(n819) );
  XOR2X1 U876 ( .IN1(n870), .IN2(N309), .Q(n869) );
  AO22X1 U877 ( .IN1(N29), .IN2(n780), .IN3(N35), .IN4(n839), .Q(n870) );
  XNOR2X1 U878 ( .IN1(keyinput23), .IN2(N11), .Q(n868) );
  XNOR2X1 U879 ( .IN1(n871), .IN2(n664), .Q(n867) );
  AO22X1 U880 ( .IN1(N29), .IN2(n690), .IN3(N27), .IN4(n839), .Q(n871) );
  MUX21X1 U881 ( .IN1(n872), .IN2(n873), .S(N29), .Q(n818) );
  NAND2X0 U882 ( .IN1(n874), .IN2(n875), .QN(n873) );
  XNOR2X1 U883 ( .IN1(n768), .IN2(N297), .Q(n875) );
  AOI221X1 U884 ( .IN1(N115), .IN2(n759), .IN3(N127), .IN4(n761), .IN5(n876), 
        .QN(n768) );
  AO22X1 U885 ( .IN1(N103), .IN2(n758), .IN3(N139), .IN4(n764), .Q(n876) );
  XNOR2X1 U886 ( .IN1(N294), .IN2(n620), .Q(n874) );
  INVX0 U887 ( .INP(n772), .ZN(n620) );
  AO221X1 U888 ( .IN1(N140), .IN2(n764), .IN3(N128), .IN4(n761), .IN5(n877), 
        .Q(n772) );
  NAND2X0 U889 ( .IN1(n878), .IN2(n879), .QN(n877) );
  XNOR2X1 U890 ( .IN1(n880), .IN2(keyinput36), .Q(n879) );
  NAND2X0 U891 ( .IN1(N104), .IN2(n758), .QN(n880) );
  NOR2X0 U892 ( .IN1(n881), .IN2(N322), .QN(n758) );
  XOR2X1 U893 ( .IN1(n882), .IN2(keyinput17), .Q(n878) );
  NAND2X0 U894 ( .IN1(N116), .IN2(n759), .QN(n882) );
  NOR2X0 U895 ( .IN1(N319), .IN2(N322), .QN(n764) );
  NAND3X0 U896 ( .IN1(n883), .IN2(n884), .IN3(n840), .QN(n872) );
  AND2X1 U897 ( .IN1(N28), .IN2(n839), .Q(n840) );
  XNOR2X1 U898 ( .IN1(N29), .IN2(keyinput21), .Q(n839) );
  XNOR2X1 U899 ( .IN1(N33), .IN2(n603), .Q(n884) );
  INVX0 U900 ( .INP(N297), .ZN(n603) );
  XNOR2X1 U901 ( .IN1(n598), .IN2(N26), .Q(n883) );
  MUX21X1 U902 ( .IN1(n885), .IN2(n886), .S(n834), .Q(n817) );
  INVX0 U903 ( .INP(N16), .ZN(n834) );
  NAND3X0 U904 ( .IN1(n887), .IN2(n888), .IN3(n889), .QN(n886) );
  XNOR2X1 U905 ( .IN1(N4), .IN2(n601), .Q(n889) );
  XNOR2X1 U906 ( .IN1(N5), .IN2(n665), .Q(n888) );
  INVX0 U907 ( .INP(N266), .ZN(n665) );
  XOR2X1 U908 ( .IN1(N256), .IN2(N19), .Q(n887) );
  NAND3X0 U909 ( .IN1(n890), .IN2(n891), .IN3(n892), .QN(n885) );
  XNOR2X1 U910 ( .IN1(n591), .IN2(N256), .Q(n892) );
  XNOR2X1 U911 ( .IN1(N1821), .IN2(N266), .Q(n891) );
  XNOR2X1 U912 ( .IN1(n596), .IN2(N259), .Q(n890) );
  XOR3X1 U913 ( .IN1(keyinput86), .IN2(n893), .IN3(n894), .Q(N2970) );
  XNOR2X1 U914 ( .IN1(N313), .IN2(n895), .Q(n894) );
  OA21X1 U915 ( .IN1(n896), .IN2(n897), .IN3(n898), .Q(n895) );
  XOR2X1 U916 ( .IN1(keyinput64), .IN2(n899), .Q(n898) );
  NOR2X0 U917 ( .IN1(n900), .IN2(n901), .QN(n899) );
  XNOR2X1 U918 ( .IN1(n902), .IN2(n903), .Q(n901) );
  INVX0 U919 ( .INP(n897), .ZN(n900) );
  AO21X1 U920 ( .IN1(N297), .IN2(n664), .IN3(n904), .Q(n897) );
  XOR2X1 U921 ( .IN1(keyinput25), .IN2(n905), .Q(n904) );
  NOR2X0 U922 ( .IN1(n906), .IN2(n664), .QN(n905) );
  XNOR2X1 U923 ( .IN1(N297), .IN2(keyinput19), .Q(n906) );
  INVX0 U924 ( .INP(N301), .ZN(n664) );
  XOR2X1 U925 ( .IN1(n902), .IN2(n903), .Q(n896) );
  AOI21X1 U926 ( .IN1(N309), .IN2(n907), .IN3(n908), .QN(n903) );
  XOR2X1 U927 ( .IN1(keyinput26), .IN2(n909), .Q(n908) );
  NOR2X0 U928 ( .IN1(n910), .IN2(n907), .QN(n909) );
  XNOR2X1 U929 ( .IN1(N309), .IN2(keyinput20), .Q(n910) );
  INVX0 U930 ( .INP(N305), .ZN(n907) );
  AO21X1 U931 ( .IN1(N355), .IN2(n598), .IN3(n911), .Q(n902) );
  XOR2X1 U932 ( .IN1(keyinput18), .IN2(n912), .Q(n911) );
  NOR2X0 U933 ( .IN1(n598), .IN2(n913), .QN(n912) );
  XOR2X1 U934 ( .IN1(keyinput7), .IN2(N355), .Q(n913) );
  INVX0 U935 ( .INP(N294), .ZN(n598) );
  AND2X1 U936 ( .IN1(N14), .IN2(n914), .Q(N2925) );
  XOR2X1 U937 ( .IN1(n915), .IN2(n916), .Q(n914) );
  MUX41X1 U938 ( .IN1(n917), .IN3(n918), .IN2(n918), .IN4(n917), .S0(N349), 
        .S1(N346), .Q(n916) );
  XOR2X1 U939 ( .IN1(n917), .IN2(keyinput45), .Q(n918) );
  AOI21X1 U940 ( .IN1(N256), .IN2(n601), .IN3(n919), .QN(n917) );
  XOR2X1 U941 ( .IN1(keyinput27), .IN2(n920), .Q(n919) );
  NOR2X0 U942 ( .IN1(N256), .IN2(n601), .QN(n920) );
  INVX0 U943 ( .INP(N259), .ZN(n601) );
  NAND3X0 U944 ( .IN1(n921), .IN2(n922), .IN3(n923), .QN(n915) );
  MUX21X1 U945 ( .IN1(n924), .IN2(n925), .S(n926), .Q(n923) );
  NAND2X0 U946 ( .IN1(n927), .IN2(n928), .QN(n925) );
  NOR2X0 U947 ( .IN1(keyinput43), .IN2(n929), .QN(n924) );
  XOR2X1 U948 ( .IN1(n930), .IN2(n931), .Q(n929) );
  OR2X1 U949 ( .IN1(keyinput33), .IN2(n932), .Q(n930) );
  OR2X1 U950 ( .IN1(n928), .IN2(n927), .Q(n922) );
  NOR2X0 U951 ( .IN1(n931), .IN2(n932), .QN(n927) );
  INVX0 U952 ( .INP(keyinput43), .ZN(n928) );
  XOR2X1 U953 ( .IN1(n933), .IN2(keyinput44), .Q(n921) );
  NAND3X0 U954 ( .IN1(n932), .IN2(n926), .IN3(n934), .QN(n933) );
  XOR2X1 U955 ( .IN1(n931), .IN2(keyinput33), .Q(n934) );
  XOR2X1 U956 ( .IN1(n935), .IN2(N331), .Q(n931) );
  NAND2X0 U957 ( .IN1(keyinput5), .IN2(N328), .QN(n935) );
  XNOR2X1 U958 ( .IN1(n936), .IN2(N343), .Q(n926) );
  NAND2X0 U959 ( .IN1(keyinput6), .IN2(N340), .QN(n936) );
  AOI21X1 U960 ( .IN1(N337), .IN2(n937), .IN3(n938), .QN(n932) );
  XOR2X1 U961 ( .IN1(n939), .IN2(keyinput10), .Q(n938) );
  OR2X1 U962 ( .IN1(n937), .IN2(N337), .Q(n939) );
  INVX0 U963 ( .INP(N334), .ZN(n937) );
  AO221X1 U964 ( .IN1(keyinput84), .IN2(n940), .IN3(n941), .IN4(n757), .IN5(
        n942), .Q(N2891) );
  XOR2X1 U965 ( .IN1(keyinput59), .IN2(n943), .Q(n942) );
  AND2X1 U966 ( .IN1(n893), .IN2(n941), .Q(n943) );
  XOR2X1 U967 ( .IN1(n944), .IN2(keyinput49), .Q(n941) );
  NAND2X0 U968 ( .IN1(n757), .IN2(n893), .QN(n944) );
  INVX0 U969 ( .INP(N316), .ZN(n893) );
  XNOR2X1 U970 ( .IN1(n945), .IN2(keyinput41), .Q(n757) );
  NAND2X0 U971 ( .IN1(n946), .IN2(n947), .QN(n945) );
  XNOR2X1 U972 ( .IN1(N313), .IN2(n775), .Q(n940) );
  AO221X1 U973 ( .IN1(N99), .IN2(n948), .IN3(N135), .IN4(n949), .IN5(n950), 
        .Q(n775) );
  AO22X1 U974 ( .IN1(N123), .IN2(n761), .IN3(N111), .IN4(n759), .Q(n950) );
  MUX21X1 U975 ( .IN1(n688), .IN2(n747), .S(N246), .Q(N2643) );
  INVX0 U976 ( .INP(n746), .ZN(n747) );
  OAI21X1 U977 ( .IN1(n746), .IN2(N241), .IN3(n596), .QN(N2496) );
  INVX0 U978 ( .INP(n589), .ZN(n596) );
  NOR2X0 U979 ( .IN1(N230), .IN2(n589), .QN(n746) );
  MUX21X1 U980 ( .IN1(N2010), .IN2(N2014), .S(N246), .Q(N2389) );
  MUX21X1 U981 ( .IN1(n589), .IN2(N2012), .S(N246), .Q(N2387) );
  AO221X1 U982 ( .IN1(N79), .IN2(n812), .IN3(N66), .IN4(n813), .IN5(n951), .Q(
        n589) );
  AO22X1 U983 ( .IN1(N54), .IN2(n815), .IN3(N92), .IN4(n816), .Q(n951) );
  XNOR2X1 U984 ( .IN1(n952), .IN2(keyinput40), .Q(N2018) );
  NAND4X0 U985 ( .IN1(n953), .IN2(n954), .IN3(n955), .IN4(n956), .QN(n952) );
  NAND2X0 U986 ( .IN1(N87), .IN2(n957), .QN(n955) );
  NAND2X0 U987 ( .IN1(N74), .IN2(n812), .QN(n954) );
  XNOR2X1 U988 ( .IN1(n958), .IN2(keyinput30), .Q(n953) );
  NAND2X0 U989 ( .IN1(N49), .IN2(n815), .QN(n958) );
  XOR2X1 U990 ( .IN1(n959), .IN2(keyinput48), .Q(N1971) );
  AO21X1 U991 ( .IN1(N3), .IN2(N1), .IN3(n960), .Q(n959) );
  NAND2X0 U992 ( .IN1(N36), .IN2(n961), .QN(N1970) );
  INVX0 U993 ( .INP(n960), .ZN(n961) );
  NAND3X0 U994 ( .IN1(N1726), .IN2(N237), .IN3(N224), .QN(n960) );
  NAND2X0 U995 ( .IN1(N241), .IN2(n591), .QN(N1969) );
  INVX0 U996 ( .INP(n688), .ZN(n591) );
  AO221X1 U997 ( .IN1(N68), .IN2(n812), .IN3(N56), .IN4(n813), .IN5(n962), .Q(
        n688) );
  AO22X1 U998 ( .IN1(N43), .IN2(n815), .IN3(N81), .IN4(n816), .Q(n962) );
  INVX0 U999 ( .INP(N2012), .ZN(N1821) );
  INVX0 U1000 ( .INP(N2014), .ZN(N1820) );
  INVX0 U1001 ( .INP(N2016), .ZN(N1819) );
  INVX0 U1002 ( .INP(n690), .ZN(N1818) );
  AO221X1 U1003 ( .IN1(N102), .IN2(n948), .IN3(N138), .IN4(n949), .IN5(n963), 
        .Q(n690) );
  AO22X1 U1004 ( .IN1(N126), .IN2(n761), .IN3(N114), .IN4(n759), .Q(n963) );
  INVX0 U1005 ( .INP(n780), .ZN(N1817) );
  AO221X1 U1006 ( .IN1(N100), .IN2(n948), .IN3(N136), .IN4(n949), .IN5(n964), 
        .Q(n780) );
  AO22X1 U1007 ( .IN1(N124), .IN2(n761), .IN3(N112), .IN4(n759), .Q(n964) );
  INVX0 U1008 ( .INP(n777), .ZN(N1816) );
  AO221X1 U1009 ( .IN1(N137), .IN2(n949), .IN3(N113), .IN4(n759), .IN5(n965), 
        .Q(n777) );
  AO21X1 U1010 ( .IN1(N125), .IN2(n761), .IN3(n966), .Q(n965) );
  XNOR2X1 U1011 ( .IN1(n967), .IN2(keyinput32), .Q(n966) );
  NAND2X0 U1012 ( .IN1(N101), .IN2(n948), .QN(n967) );
  NOR2X0 U1013 ( .IN1(n881), .IN2(n946), .QN(n948) );
  NOR2X0 U1014 ( .IN1(n947), .IN2(N319), .QN(n761) );
  NOR2X0 U1015 ( .IN1(n881), .IN2(n947), .QN(n759) );
  INVX0 U1016 ( .INP(N319), .ZN(n881) );
  NOR2X0 U1017 ( .IN1(n946), .IN2(N319), .QN(n949) );
  XOR2X1 U1018 ( .IN1(n947), .IN2(keyinput15), .Q(n946) );
  INVX0 U1019 ( .INP(N322), .ZN(n947) );
  XNOR2X1 U1020 ( .IN1(keyinput39), .IN2(n968), .Q(N1726) );
  OA22X1 U1021 ( .IN1(n969), .IN2(n970), .IN3(n971), .IN4(n972), .Q(n968) );
  INVX0 U1022 ( .INP(N325), .ZN(n972) );
  INVX0 U1023 ( .INP(N231), .ZN(n970) );
  XOR2X1 U1024 ( .IN1(n973), .IN2(keyinput11), .Q(n969) );
  AO221X1 U1025 ( .IN1(N85), .IN2(n974), .IN3(N60), .IN4(n975), .IN5(n976), 
        .Q(N2022) );
  AO21X1 U1026 ( .IN1(N72), .IN2(n812), .IN3(n977), .Q(n976) );
  XNOR2X1 U1027 ( .IN1(n978), .IN2(keyinput31), .Q(n977) );
  NAND2X0 U1028 ( .IN1(N47), .IN2(n815), .QN(n978) );
  AO221X1 U1029 ( .IN1(N86), .IN2(n974), .IN3(N61), .IN4(n975), .IN5(n979), 
        .Q(N2020) );
  AO22X1 U1030 ( .IN1(N73), .IN2(n812), .IN3(N48), .IN4(n815), .Q(n979) );
  AO221X1 U1031 ( .IN1(N88), .IN2(n974), .IN3(N62), .IN4(n975), .IN5(n980), 
        .Q(N2016) );
  AO22X1 U1032 ( .IN1(N75), .IN2(n812), .IN3(N50), .IN4(n815), .Q(n980) );
  AO221X1 U1033 ( .IN1(N89), .IN2(n974), .IN3(N63), .IN4(n975), .IN5(n981), 
        .Q(N2014) );
  AO21X1 U1034 ( .IN1(N51), .IN2(n815), .IN3(n982), .Q(n981) );
  XOR2X1 U1035 ( .IN1(n983), .IN2(keyinput14), .Q(n982) );
  NAND2X0 U1036 ( .IN1(N76), .IN2(n812), .QN(n983) );
  INVX0 U1037 ( .INP(n956), .ZN(n975) );
  NAND2X0 U1038 ( .IN1(N234), .IN2(n957), .QN(n956) );
  AND2X1 U1039 ( .IN1(n957), .IN2(n984), .Q(n974) );
  XNOR2X1 U1040 ( .IN1(n985), .IN2(keyinput13), .Q(n957) );
  AO221X1 U1041 ( .IN1(N77), .IN2(n812), .IN3(N64), .IN4(n813), .IN5(n986), 
        .Q(N2012) );
  AO22X1 U1042 ( .IN1(N52), .IN2(n815), .IN3(N90), .IN4(n816), .Q(n986) );
  AO221X1 U1043 ( .IN1(N53), .IN2(n815), .IN3(N78), .IN4(n812), .IN5(n987), 
        .Q(N2010) );
  AO21X1 U1044 ( .IN1(N65), .IN2(n813), .IN3(n988), .Q(n987) );
  XOR2X1 U1045 ( .IN1(n989), .IN2(keyinput29), .Q(n988) );
  NAND2X0 U1046 ( .IN1(N91), .IN2(n816), .QN(n989) );
  MUX21X1 U1047 ( .IN1(n815), .IN2(n990), .S(keyinput12), .Q(n816) );
  NOR2X0 U1048 ( .IN1(N227), .IN2(N234), .QN(n990) );
  MUX21X1 U1049 ( .IN1(n812), .IN2(n991), .S(keyinput12), .Q(n813) );
  NOR2X0 U1050 ( .IN1(n984), .IN2(N227), .QN(n991) );
  NOR2X0 U1051 ( .IN1(n984), .IN2(n985), .QN(n812) );
  INVX0 U1052 ( .INP(N234), .ZN(n984) );
  NOR2X0 U1053 ( .IN1(n985), .IN2(N234), .QN(n815) );
  INVX0 U1054 ( .INP(N227), .ZN(n985) );
  INVX0 U1055 ( .INP(N1448), .ZN(N1277) );
  NAND2X0 U1056 ( .IN1(n971), .IN2(n973), .QN(N1448) );
  XOR2X1 U1057 ( .IN1(n992), .IN2(keyinput4), .Q(n973) );
  NAND4X0 U1058 ( .IN1(N57), .IN2(N69), .IN3(N120), .IN4(N108), .QN(n992) );
  AND4X1 U1059 ( .IN1(N44), .IN2(N132), .IN3(N82), .IN4(N96), .Q(n971) );
  XOR2X1 U1060 ( .IN1(n993), .IN2(keyinput22), .Q(N1269) );
  NAND2X0 U1061 ( .IN1(N325), .IN2(n994), .QN(n993) );
  NAND2X0 U1062 ( .IN1(N231), .IN2(n994), .QN(N1029) );
  INVX0 U1063 ( .INP(N1028), .ZN(n994) );
  NAND2X0 U1064 ( .IN1(N7), .IN2(N237), .QN(N1028) );
  AND2X1 U1065 ( .IN1(N94), .IN2(N219), .Q(N1026) );
endmodule

