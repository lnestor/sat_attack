// Verilog File 
module c1908_lut_128bit.bench (G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput1_7,keyinput0_7,keyinput0_2,keyinput0_4,keyinput0_3,keyinput0_1,
keyinput0_5,keyinput0_0,keyinput1_0,keyinput2_0,keyinput3_0,keyinput4_0,keyinput5_0,keyinput6_0,keyinput7_0,keyinput8_0,
keyinput9_0,keyinput10_0,keyinput11_0,keyinput12_0,keyinput13_0,keyinput14_0,keyinput15_0,keyinput1_1,keyinput2_1,keyinput3_1,
keyinput4_1,keyinput5_1,keyinput6_1,keyinput7_1,keyinput8_1,keyinput9_1,keyinput10_1,keyinput11_1,keyinput12_1,keyinput13_1,
keyinput14_1,keyinput15_1,keyinput1_2,keyinput2_2,keyinput3_2,keyinput4_2,keyinput5_2,keyinput6_2,keyinput7_2,keyinput8_2,
keyinput9_2,keyinput10_2,keyinput11_2,keyinput12_2,keyinput13_2,keyinput14_2,keyinput15_2,keyinput1_3,keyinput2_3,keyinput3_3,
keyinput4_3,keyinput5_3,keyinput6_3,keyinput7_3,keyinput8_3,keyinput9_3,keyinput10_3,keyinput11_3,keyinput12_3,keyinput13_3,
keyinput14_3,keyinput15_3,keyinput1_4,keyinput2_4,keyinput3_4,keyinput4_4,keyinput5_4,keyinput6_4,keyinput7_4,keyinput8_4,
keyinput9_4,keyinput10_4,keyinput11_4,keyinput12_4,keyinput13_4,keyinput14_4,keyinput15_4,keyinput1_5,keyinput2_5,keyinput3_5,
keyinput4_5,keyinput5_5,keyinput6_5,keyinput7_5,keyinput8_5,keyinput9_5,keyinput10_5,keyinput11_5,keyinput12_5,keyinput13_5,
keyinput14_5,keyinput15_5,keyinput0_6,keyinput1_6,keyinput2_6,keyinput3_6,keyinput4_6,keyinput5_6,keyinput6_6,keyinput7_6,
keyinput8_6,keyinput9_6,keyinput10_6,keyinput11_6,keyinput12_6,keyinput13_6,keyinput14_6,keyinput15_6,keyinput2_7,keyinput3_7,
keyinput4_7,keyinput5_7,keyinput6_7,keyinput7_7,keyinput8_7,keyinput9_7,keyinput10_7,keyinput11_7,keyinput12_7,keyinput13_7,
keyinput14_7,keyinput15_7,G3,G6,G9,G12,G30,G45,G48,G15,
G18,G21,G24,G27,G33,G36,G39,G42,G75,G51,
G54,G60,G63,G66,G69,G72,G57);

input G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,keyinput1_7,keyinput0_7,keyinput0_2,keyinput0_4,keyinput0_3,keyinput0_1,
keyinput0_5,keyinput0_0,keyinput1_0,keyinput2_0,keyinput3_0,keyinput4_0,keyinput5_0,keyinput6_0,keyinput7_0,keyinput8_0,
keyinput9_0,keyinput10_0,keyinput11_0,keyinput12_0,keyinput13_0,keyinput14_0,keyinput15_0,keyinput1_1,keyinput2_1,keyinput3_1,
keyinput4_1,keyinput5_1,keyinput6_1,keyinput7_1,keyinput8_1,keyinput9_1,keyinput10_1,keyinput11_1,keyinput12_1,keyinput13_1,
keyinput14_1,keyinput15_1,keyinput1_2,keyinput2_2,keyinput3_2,keyinput4_2,keyinput5_2,keyinput6_2,keyinput7_2,keyinput8_2,
keyinput9_2,keyinput10_2,keyinput11_2,keyinput12_2,keyinput13_2,keyinput14_2,keyinput15_2,keyinput1_3,keyinput2_3,keyinput3_3,
keyinput4_3,keyinput5_3,keyinput6_3,keyinput7_3,keyinput8_3,keyinput9_3,keyinput10_3,keyinput11_3,keyinput12_3,keyinput13_3,
keyinput14_3,keyinput15_3,keyinput1_4,keyinput2_4,keyinput3_4,keyinput4_4,keyinput5_4,keyinput6_4,keyinput7_4,keyinput8_4,
keyinput9_4,keyinput10_4,keyinput11_4,keyinput12_4,keyinput13_4,keyinput14_4,keyinput15_4,keyinput1_5,keyinput2_5,keyinput3_5,
keyinput4_5,keyinput5_5,keyinput6_5,keyinput7_5,keyinput8_5,keyinput9_5,keyinput10_5,keyinput11_5,keyinput12_5,keyinput13_5,
keyinput14_5,keyinput15_5,keyinput0_6,keyinput1_6,keyinput2_6,keyinput3_6,keyinput4_6,keyinput5_6,keyinput6_6,keyinput7_6,
keyinput8_6,keyinput9_6,keyinput10_6,keyinput11_6,keyinput12_6,keyinput13_6,keyinput14_6,keyinput15_6,keyinput2_7,keyinput3_7,
keyinput4_7,keyinput5_7,keyinput6_7,keyinput7_7,keyinput8_7,keyinput9_7,keyinput10_7,keyinput11_7,keyinput12_7,keyinput13_7,
keyinput14_7,keyinput15_7;


output G3, G6, G9, G12, G30, G45, G48, G15, G18, 
G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, 
G60, G63, G66, G69, G72, G57;

wire G149, G153, G156, G160, G165, G168, G171, G175, G179, 
G184, G188, G191, G194, G198, G202, G206, G231, G233, G241, 
G244, G245, G248, G517, G529, G541, G553, G859, G862, G907, 
G909, G911, G918, G919, G922, G926, G930, G932, G934, G938, 
G943, G947, G949, G1506, G1514, G1522, G1530, G1538, G1546, G1554, 
G1562, G1570, G1578, G1586, G1594, G1602, G1610, G1618, G1626, G1512, 
G1520, G1528, G1536, G1544, G1552, G1560, G1568, G1576, G1584, G1592, 
G1600, G1608, G1616, G1624, G1632, G50, G52, G56, G58, G62, 
G64, G251, G254, G288, G291, G299, G302, G318, G321, G327, 
G330, G352, G355, G369, G382, G385, G853, G856, G893, G954, 
G955, G1050, G1053, G1176, G1179, G1197, G1207, G1222, G1244, G1278, 
G1290, G1300, G1312, G1332, G1335, G1442, G1450, G1458, G1466, G1474, 
G1482, G1490, G1498, G1634, G1644, G1657, G1665, G1697, G1705, G1713, 
G1721, G1745, G1753, G1785, G1793, G1814, G1817, G1830, G1833, G1841, 
G1849, G1854, G1857, G1870, G1873, G1878, G1881, G1642, G1652, G1056, 
G1057, G1182, G1183, G1211, G1298, G1320, G1338, G1339, G457, G459, 
G482, G487, G492, G505, G1456, G1448, G1472, G1464, G1488, G1480, 
G1504, G1496, G967, G978, G979, G980, G1661, G990, G1669, G1030, 
G1701, G1040, G1709, G1058, G1717, G1068, G1725, G1078, G1090, G1100, 
G1749, G1112, G1757, G1154, G1789, G1166, G1797, G1194, G1201, G1204, 
G1820, G1821, G1230, G1836, G1837, G1252, G1256, G1845, G1268, G1853, 
G1860, G1861, G1286, G1876, G1877, G1308, G1884, G1885, G1654, G1662, 
G1694, G1702, G1710, G1718, G1726, G1734, G1742, G1750, G1782, G1790, 
G1838, G1846, G297, G298, G361, G362, G404, G405, G1225, G1226, 
G1247, G1248, G1281, G1282, G1303, G1304, G998, G988, G268, G1038, 
G1048, G1076, G1066, G1098, G1120, G1174, G363, G1210, G373, G1276, 
G406, G565, G566, G614, G615, G956, G958, G969, G1660, G984, 
G1668, G994, G1700, G1034, G1708, G1044, G1716, G1062, G1724, G1072, 
G1732, G1086, G1740, G1748, G1104, G1108, G1756, G1116, G1788, G1158, 
G1162, G1796, G1170, G1200, G1203, G1227, G1249, G1844, G1260, G1264, 
G1852, G1272, G1283, G1305, G1410, G1418, G1426, G1434, G269, G372, 
G983, G993, G1033, G1043, G1061, G1071, G1103, G1115, G1157, G1169, 
G1184, G1202, G1259, G1271, G1322, G374, G1317, G396, G1321, G1424, 
G1416, G1440, G1432, G985, G995, G1035, G1045, G1063, G1073, G1105, 
G1117, G1159, G1171, G1212, G1231, G1232, G1253, G1254, G1261, G1273, 
G1287, G1288, G1309, G1310, G1192, G397, G1330, G1000, G1010, G1233, 
G1255, G1289, G1311, G1381, G257, G999, G989, G272, G1039, G294, 
G1049, G305, G1077, G308, G1067, G1121, G358, G1175, G1220, G388, 
G1277, G398, G1109, G1110, G1163, G1164, G1234, G1265, G1266, G1822, 
G1862, G1865, G258, G273, G1018, G1008, G295, G306, G309, G359, 
G389, G1385, G1111, G1165, G1267, G1886, G259, G274, G296, G307, 
G310, G360, G1242, G390, G1828, G1868, G1869, G1373, G1798, G1825, 
G265, G314, G407, G1293, G1294, G1892, G1777, G1889, G410, G1377, 
G1804, G1237, G1829, G1295, G1670, G1678, G1729, G1737, G262, G1761, 
G1769, G336, G340, G343, G1781, G1238, G1325, G1893, G1340, G1352, 
G1673, G1681, G1801, G1897, G1905, G391, G1299, G1676, G1684, G1081, 
G1733, G1093, G1741, G1765, G1773, G1239, G1326, G1894, G1902, G392, 
G1360, G1003, G1677, G1013, G1685, G1082, G1094, G1122, G1134, G1187, 
G1805, G1327, G1901, G1348, G1909, G1758, G1766, G377, G1243, G393, 
G1004, G1014, G1083, G1095, G1188, G1900, G1344, G1908, G1356, G1142, 
G378, G399, G1331, G1005, G1015, G1764, G1130, G1772, G1138, G1189, 
G1343, G1355, G324, G1099, G379, G400, G449, G1087, G1088, G1137, 
G1345, G1357, G1397, G277, G1019, G280, G1009, G325, G364, G1193, 
G401, G1089, G1139, G278, G281, G326, G365, G413, G1361, G1401, 
G445, G1349, G1350, G1389, G1493, G1501, G1689, G279, G282, G1143, 
G366, G414, G453, G1127, G1131, G1132, G1351, G1365, G1405, G285, 
G367, G415, G1393, G556, G1505, G559, G1497, G1693, G1133, G1477, 
G1485, G1809, G1369, G1409, G557, G560, G1362, G1378, G1429, G1437, 
G1686, G1774, G1910, G1918, G544, G1489, G547, G1481, G558, G561, 
G1813, G348, G1370, G1368, G1384, G424, G508, G1441, G511, G1433, 
G545, G548, G564, G1692, G1024, G1780, G1148, G1916, G1924, G1376, 
G421, G423, G509, G512, G546, G549, G719, G722, G1023, G1147, 
G420, G425, G510, G513, G552, G1025, G1149, G418, G419, G422, 
G441, G516, G725, G728, G1029, G1153, G433, G437, G663, G666, 
G731, G746, G756, G770, G1461, G1469, G1413, G1421, G1445, G1453, 
G532, G1473, G535, G1465, G495, G1425, G498, G1417, G1457, G523, 
G1449, G533, G536, G496, G499, G524, G534, G537, G497, G500, 
G525, G540, G503, G522, G528, G669, G672, G569, G588, G618, 
G639, G867, G588a, G588b, G639a, G639b, G675, G688, G696, G710, 
G73, G572, G573, G621, G622, G776, G780, G784, G788, G812, 
G832, G836, G1509, G1517, G1525, G1533, G1581, G1621, G1629, G792, 
G796, G800, G804, G808, G816, G820, G824, G828, G871, G873, 
G875, G877, G879, G881, G883, G885, G1541, G1549, G1557, G1565, 
G1573, G1589, G1597, G1605, G1613, G1, G1513, G4, G1521, G7, 
G1529, G10, G1537, G28, G1585, G43, G1625, G46, G1633, G886, 
G2, G5, G8, G11, G13, G1545, G16, G1553, G19, G1561, 
G22, G1569, G25, G1577, G29, G31, G1593, G34, G1601, G37, 
G1609, G40, G1617, G44, G47, G857, G860, G863, G865, G14, 
G17, G20, G23, G26, G32, G35, G38, G41, G1913, G1921, 
G887, G462, G74, G1637, G1917, G1647, G1925, G1020, G1144, G1386, 
G1394, G1402, G1638, G1648, G1806, G1639, G1649, G287, G350, G427, 
G429, G431, G1028, G1152, G1392, G1400, G1408, G1812, G1216, G286, 
G349, G426, G428, G430, G67, G1643, G70, G1653, G1215, G49, 
G53, G59, G61, G65, G68, G71, G1217, G375, G1221, G376, 
G55, in0not_0, in1not_0, in2not_0, in3not_0, T0_0, T1_0, T2_0, T3_0, T4_0, 
T5_0, T6_0, T7_0, T8_0, T9_0, T10_0, T11_0, T12_0, T13_0, T14_0, 
T15_0, in0not_1, in1not_1, in2not_1, in3not_1, T0_1, T1_1, T2_1, T3_1, T4_1, 
T5_1, T6_1, T7_1, T8_1, T9_1, T10_1, T11_1, T12_1, T13_1, T14_1, 
T15_1, in0not_2, in1not_2, in2not_2, in3not_2, T0_2, T1_2, T2_2, T3_2, T4_2, 
T5_2, T6_2, T7_2, T8_2, T9_2, T10_2, T11_2, T12_2, T13_2, T14_2, 
T15_2, in0not_3, in1not_3, in2not_3, in3not_3, T0_3, T1_3, T2_3, T3_3, T4_3, 
T5_3, T6_3, T7_3, T8_3, T9_3, T10_3, T11_3, T12_3, T13_3, T14_3, 
T15_3, in0not_4, in1not_4, in2not_4, in3not_4, T0_4, T1_4, T2_4, T3_4, T4_4, 
T5_4, T6_4, T7_4, T8_4, T9_4, T10_4, T11_4, T12_4, T13_4, T14_4, 
T15_4, in0not_5, in1not_5, in2not_5, in3not_5, T0_5, T1_5, T2_5, T3_5, T4_5, 
T5_5, T6_5, T7_5, T8_5, T9_5, T10_5, T11_5, T12_5, T13_5, T14_5, 
T15_5, in0not_6, in1not_6, in2not_6, in3not_6, T0_6, T1_6, T2_6, T3_6, T4_6, 
T5_6, T6_6, T7_6, T8_6, T9_6, T10_6, T11_6, T12_6, T13_6, T14_6, 
T15_6, in0not_7, in1not_7, in2not_7, in3not_7, T0_7, T1_7, T2_7, T3_7, T4_7, 
T5_7, T6_7, T7_7, T8_7, T9_7, T10_7, T11_7, T12_7, T13_7, T14_7, 
T15_7;

not g0(G149, G101);
not g1(G153, G104);
not g2(G156, G107);
not g3(G160, G110);
not g4(G165, G113);
not g5(G168, G116);
not g6(G171, G119);
not g7(G175, G122);
not g8(G179, G125);
not g9(G184, G128);
not g10(G188, G131);
not g11(G191, G134);
not g12(G194, G137);
not g13(G198, G140);
not g14(G202, G143);
not g15(G206, G146);
nand g16(G231, G224, G898);
nand g17(G233, G227, G900);
not g18(G241, G237);
not g19(G244, G237);
assign G245 = G234;
assign G248 = G234;
not g22(G517, G469);
not g23(G529, G472);
not g24(G541, G475);
not g25(G553, G478);
not g26(G859, G953);
not g27(G862, G953);
not g28(G907, G898);
not g29(G909, G900);
assign G911 = G902;
not g31(G918, G902);
assign G919 = G902;
not g33(G922, G902);
assign G926 = G952;
not g35(G930, G952);
not g36(G932, G952);
assign G934 = G953;
not g38(G938, G953);
assign G943 = G953;
assign G947 = G953;
not g41(G949, G953);
assign G1506 = G101;
assign G1514 = G104;
assign G1522 = G107;
assign G1530 = G110;
assign G1538 = G113;
assign G1546 = G116;
assign G1554 = G119;
assign G1562 = G122;
assign G1570 = G125;
assign G1578 = G128;
assign G1586 = G131;
assign G1594 = G134;
assign G1602 = G137;
assign G1610 = G140;
assign G1618 = G143;
assign G1626 = G146;
not g58(G1512, G1506);
not g59(G1520, G1514);
not g60(G1528, G1522);
not g61(G1536, G1530);
not g62(G1544, G1538);
not g63(G1552, G1546);
not g64(G1560, G1554);
not g65(G1568, G1562);
not g66(G1576, G1570);
not g67(G1584, G1578);
not g68(G1592, G1586);
not g69(G1600, G1594);
not g70(G1608, G1602);
not g71(G1616, G1610);
not g72(G1624, G1618);
not g73(G1632, G1626);
nand g74(G50, G930, G947);
nand g75(G52, G930, G947);
nand g76(G56, G930, G947);
nand g77(G58, G930, G947);
nand g78(G62, G930, G947);
nand g79(G64, G930, G947);
assign G251 = G149;
assign G254 = G153;
assign G288 = G165;
assign G291 = G168;
assign G299 = G184;
assign G302 = G202;
and g86(G318, G224, G938);
assign G321 = G179;
assign G327 = G188;
assign G330 = G191;
and g90(G352, G227, G938);
assign G355 = G198;
and g92(G369, G210, G241, G938);
assign G382 = G206;
assign G385 = G198;
nand g95(G853, G943, G907);
nand g96(G856, G943, G909);
nand g97(G893, G248, G237);
nand g98(G954, G248, G922);
nand g99(G955, G244, G922);
assign G1050 = G160;
assign G1053 = G175;
assign G1176 = G179;
assign G1179 = G198;
assign G1197 = G149;
assign G1207 = G149;
assign G1222 = G153;
assign G1244 = G188;
assign G1278 = G156;
and g109(G1290, G217, G245, G938);
assign G1300 = G191;
assign G1312 = G160;
assign G1332 = G194;
and g113(G1335, G221, G245, G938);
assign G1442 = G517;
assign G1450 = G517;
assign G1458 = G529;
assign G1466 = G529;
assign G1474 = G541;
assign G1482 = G541;
assign G1490 = G553;
assign G1498 = G553;
and g122(G1634, G231, G934);
and g123(G1644, G233, G934);
assign G1657 = G156;
assign G1665 = G156;
assign G1697 = G171;
assign G1705 = G171;
assign G1713 = G206;
assign G1721 = G206;
assign G1745 = G194;
assign G1753 = G194;
assign G1785 = G160;
assign G1793 = G160;
assign G1814 = G165;
assign G1817 = G175;
and g136(G1830, G214, G241, G938);
assign G1833 = G202;
assign G1841 = G179;
assign G1849 = G179;
assign G1854 = G168;
assign G1857 = G175;
assign G1870 = G184;
assign G1873 = G202;
assign G1878 = G171;
assign G1881 = G184;
not g146(G1642, G1634);
not g147(G1652, G1644);
not g148(G1056, G1050);
not g149(G1057, G1053);
not g150(G1182, G1176);
not g151(G1183, G1179);
not g152(G1211, G1207);
not g153(G1298, G1290);
not g154(G1320, G1312);
not g155(G1338, G1332);
not g156(G1339, G1335);
and g157(G457, G210, G955);
and g158(G459, G217, G954);
nand g159(G482, G214, G955);
nand g160(G487, G221, G954);
nand g161(G492, G210, G955);
nand g162(G505, G217, G954);
not g163(G1456, G1450);
not g164(G1448, G1442);
not g165(G1472, G1466);
not g166(G1464, G1458);
not g167(G1488, G1482);
not g168(G1480, G1474);
not g169(G1504, G1498);
not g170(G1496, G1490);
nand g171(G967, G909, G919, G943, G893);
nand g172(G978, G926, G949, G893);
and g173(G979, G926, G949, G893);
assign G980 = G251;
not g175(G1661, G1657);
assign G990 = G251;
not g177(G1669, G1665);
assign G1030 = G288;
not g179(G1701, G1697);
assign G1040 = G288;
not g181(G1709, G1705);
assign G1058 = G299;
not g183(G1717, G1713);
assign G1068 = G299;
not g185(G1725, G1721);
assign G1078 = G318;
assign G1090 = G318;
assign G1100 = G327;
not g189(G1749, G1745);
assign G1112 = G327;
not g191(G1757, G1753);
assign G1154 = G352;
not g193(G1789, G1785);
assign G1166 = G352;
not g195(G1797, G1793);
assign G1194 = G369;
not g197(G1201, G1197);
assign G1204 = G369;
not g199(G1820, G1814);
not g200(G1821, G1817);
not g201(G1230, G1222);
not g202(G1836, G1830);
not g203(G1837, G1833);
not g204(G1252, G1244);
assign G1256 = G382;
not g206(G1845, G1841);
assign G1268 = G382;
not g208(G1853, G1849);
not g209(G1860, G1854);
not g210(G1861, G1857);
not g211(G1286, G1278);
not g212(G1876, G1870);
not g213(G1877, G1873);
not g214(G1308, G1300);
not g215(G1884, G1878);
not g216(G1885, G1881);
assign G1654 = G254;
assign G1662 = G254;
assign G1694 = G291;
assign G1702 = G291;
assign G1710 = G302;
assign G1718 = G302;
assign G1726 = G321;
assign G1734 = G321;
assign G1742 = G330;
assign G1750 = G330;
assign G1782 = G355;
assign G1790 = G355;
assign G1838 = G385;
assign G1846 = G385;
nand g231(G297, G1053, G1056);
nand g232(G298, G1050, G1057);
nand g233(G361, G1179, G1182);
nand g234(G362, G1176, G1183);
nand g235(G404, G1335, G1338);
nand g236(G405, G1332, G1339);
nand g237(G1225, G1817, G1820);
nand g238(G1226, G1814, G1821);
nand g239(G1247, G1833, G1836);
nand g240(G1248, G1830, G1837);
nand g241(G1281, G1857, G1860);
nand g242(G1282, G1854, G1861);
nand g243(G1303, G1873, G1876);
nand g244(G1304, G1870, G1877);
not g245(G998, G990);
not g246(G988, G980);
nand g247(G268, G297, G298);
not g248(G1038, G1030);
not g249(G1048, G1040);
not g250(G1076, G1068);
not g251(G1066, G1058);
not g252(G1098, G1090);
not g253(G1120, G1112);
not g254(G1174, G1166);
nand g255(G363, G361, G362);
not g256(G1210, G1204);
nand g257(G373, G1204, G1211);
not g258(G1276, G1268);
nand g259(G406, G404, G405);
not g260(G565, G482);
assign G566 = G482;
not g262(G614, G487);
assign G615 = G487;
nand g264(G958, G956, G978);
nand g265(G969, G967, G978);
not g266(G1660, G1654);
nand g267(G984, G1654, G1661);
not g268(G1668, G1662);
nand g269(G994, G1662, G1669);
not g270(G1700, G1694);
nand g271(G1034, G1694, G1701);
not g272(G1708, G1702);
nand g273(G1044, G1702, G1709);
not g274(G1716, G1710);
nand g275(G1062, G1710, G1717);
not g276(G1724, G1718);
nand g277(G1072, G1718, G1725);
not g278(G1732, G1726);
not g279(G1086, G1078);
not g280(G1740, G1734);
not g281(G1748, G1742);
nand g282(G1104, G1742, G1749);
not g283(G1108, G1100);
not g284(G1756, G1750);
nand g285(G1116, G1750, G1757);
not g286(G1788, G1782);
nand g287(G1158, G1782, G1789);
not g288(G1162, G1154);
not g289(G1796, G1790);
nand g290(G1170, G1790, G1797);
not g291(G1200, G1194);
nand g292(G1203, G1194, G1201);
nand g293(G1227, G1225, G1226);
nand g294(G1249, G1247, G1248);
not g295(G1844, G1838);
nand g296(G1260, G1838, G1845);
not g297(G1264, G1256);
not g298(G1852, G1846);
nand g299(G1272, G1846, G1853);
nand g300(G1283, G1281, G1282);
nand g301(G1305, G1303, G1304);
assign G1410 = G492;
assign G1418 = G492;
assign G1426 = G505;
assign G1434 = G505;
not g306(G269, G268);
nand g307(G372, G1207, G1210);
nand g308(G983, G1657, G1660);
nand g309(G993, G1665, G1668);
nand g310(G1033, G1697, G1700);
nand g311(G1043, G1705, G1708);
nand g312(G1061, G1713, G1716);
nand g313(G1071, G1721, G1724);
nand g314(G1103, G1745, G1748);
nand g315(G1115, G1753, G1756);
nand g316(G1157, G1785, G1788);
nand g317(G1169, G1793, G1796);
not g318(G1184, G363);
nand g319(G1202, G1197, G1200);
nand g320(G1259, G1841, G1844);
nand g321(G1271, G1849, G1852);
not g322(G1322, G406);
nand g323(G374, G372, G373);
nand g324(G396, G1317, G1320);
not g325(G1321, G1317);
not g326(G1424, G1418);
not g327(G1416, G1410);
not g328(G1440, G1434);
not g329(G1432, G1426);
nand g330(G985, G983, G984);
nand g331(G995, G993, G994);
nand g332(G1035, G1033, G1034);
nand g333(G1045, G1043, G1044);
nand g334(G1063, G1061, G1062);
nand g335(G1073, G1071, G1072);
nand g336(G1105, G1103, G1104);
nand g337(G1117, G1115, G1116);
nand g338(G1159, G1157, G1158);
nand g339(G1171, G1169, G1170);
nand g340(G1212, G1202, G1203);
not g341(G1231, G1227);
nand g342(G1232, G1227, G1230);
not g343(G1253, G1249);
nand g344(G1254, G1249, G1252);
nand g345(G1261, G1259, G1260);
nand g346(G1273, G1271, G1272);
not g347(G1287, G1283);
nand g348(G1288, G1283, G1286);
not g349(G1309, G1305);
nand g350(G1310, G1305, G1308);
not g351(G1192, G1184);
nand g352(G397, G1312, G1321);
not g353(G1330, G1322);
assign G1000 = G269;
assign G1010 = G269;
nand g356(G1233, G1222, G1231);
nand g357(G1255, G1244, G1253);
nand g358(G1289, G1278, G1287);
nand g359(G1311, G1300, G1309);
not g360(G1381, G374);
nand g361(G257, G995, G998);
not g362(G999, G995);
not g363(G989, G985);
nand g364(G272, G1035, G1038);
not g365(G1039, G1035);
nand g366(G294, G1045, G1048);
not g367(G1049, G1045);
nand g368(G305, G1073, G1076);
not g369(G1077, G1073);
nand g370(G308, G1063, G1066);
not g371(G1067, G1063);
not g372(G1121, G1117);
nand g373(G358, G1171, G1174);
not g374(G1175, G1171);
not g375(G1220, G1212);
nand g376(G388, G1273, G1276);
not g377(G1277, G1273);
nand g378(G398, G396, G397);
not g379(G1109, G1105);
nand g380(G1110, G1105, G1108);
not g381(G1163, G1159);
nand g382(G1164, G1159, G1162);
nand g383(G1234, G1232, G1233);
not g384(G1265, G1261);
nand g385(G1266, G1261, G1264);
nand g386(G1822, G1254, G1255);
nand g387(G1862, G1310, G1311);
nand g388(G1865, G1288, G1289);
nand g389(G258, G990, G999);
nand g390(G273, G1030, G1039);
not g391(G1018, G1010);
not g392(G1008, G1000);
nand g393(G295, G1040, G1049);
nand g394(G306, G1068, G1077);
nand g395(G309, G1058, G1067);
nand g396(G359, G1166, G1175);
nand g397(G389, G1268, G1277);
not g398(G1385, G1381);
nand g399(G1111, G1100, G1109);
nand g400(G1165, G1154, G1163);
nand g401(G1267, G1256, G1265);
not g402(G1886, G398);
nand g403(G259, G257, G258);
nand g404(G274, G272, G273);
nand g405(G296, G294, G295);
nand g406(G307, G305, G306);
nand g407(G310, G308, G309);
nand g408(G360, G358, G359);
not g409(G1242, G1234);
nand g410(G390, G388, G389);
not g411(G1828, G1822);
not g412(G1868, G1862);
not g413(G1869, G1865);
nand g414(G1373, G1164, G1165);
nand g415(G1798, G1110, G1111);
nand g416(G1825, G1266, G1267);
not g417(G265, G259);
not g418(G314, G307);
not g419(G407, G296);
nand g420(G1293, G1865, G1868);
nand g421(G1294, G1862, G1869);
not g422(G1892, G1886);
not g423(G1777, G360);
not g424(G1889, G390);
assign G410 = G310;
not g426(G1377, G1373);
not g427(G1804, G1798);
nand g428(G1237, G1825, G1828);
not g429(G1829, G1825);
nand g430(G1295, G1293, G1294);
assign G1670 = G274;
assign G1678 = G274;
assign G1729 = G310;
assign G1737 = G310;
assign G1761 = G262;
assign G1769 = G262;
assign G340 = G336;
assign G343 = G314;
not g439(G1781, G1777);
nand g440(G1238, G1822, G1829);
nand g441(G1325, G1889, G1892);
not g442(G1893, G1889);
assign G1340 = G407;
assign G1352 = G407;
assign G1673 = G265;
assign G1681 = G265;
assign G1801 = G314;
assign G1897 = G336;
assign G1905 = G336;
nand g450(G391, G1295, G1298);
not g451(G1299, G1295);
not g452(G1676, G1670);
not g453(G1684, G1678);
nand g454(G1081, G1729, G1732);
not g455(G1733, G1729);
nand g456(G1093, G1737, G1740);
not g457(G1741, G1737);
not g458(G1765, G1761);
not g459(G1773, G1769);
nand g460(G1239, G1237, G1238);
nand g461(G1326, G1886, G1893);
assign G1894 = G410;
assign G1902 = G410;
nand g464(G392, G1290, G1299);
not g465(G1360, G1352);
nand g466(G1003, G1673, G1676);
not g467(G1677, G1673);
nand g468(G1013, G1681, G1684);
not g469(G1685, G1681);
nand g470(G1082, G1726, G1733);
nand g471(G1094, G1734, G1741);
assign G1122 = G340;
assign G1134 = G340;
nand g474(G1187, G1801, G1804);
not g475(G1805, G1801);
nand g476(G1327, G1325, G1326);
not g477(G1901, G1897);
not g478(G1348, G1340);
not g479(G1909, G1905);
assign G1758 = G343;
assign G1766 = G343;
nand g482(G377, G1239, G1242);
not g483(G1243, G1239);
nand g484(G393, G391, G392);
nand g485(G1004, G1670, G1677);
nand g486(G1014, G1678, G1685);
nand g487(G1083, G1081, G1082);
nand g488(G1095, G1093, G1094);
nand g489(G1188, G1798, G1805);
not g490(G1900, G1894);
nand g491(G1344, G1894, G1901);
not g492(G1908, G1902);
nand g493(G1356, G1902, G1909);
not g494(G1142, G1134);
nand g495(G378, G1234, G1243);
nand g496(G399, G1327, G1330);
not g497(G1331, G1327);
nand g498(G1005, G1003, G1004);
nand g499(G1015, G1013, G1014);
not g500(G1764, G1758);
not g501(G1130, G1122);
not g502(G1772, G1766);
nand g503(G1138, G1766, G1773);
nand g504(G1189, G1187, G1188);
nand g505(G1343, G1897, G1900);
nand g506(G1355, G1905, G1908);
nand g507(G324, G1095, G1098);
not g508(G1099, G1095);
nand g509(G379, G377, G378);
nand g510(G400, G1322, G1331);
nand g511(G449, G393, G918);
not g512(G1087, G1083);
nand g513(G1088, G1083, G1086);
nand g514(G1137, G1769, G1772);
nand g515(G1345, G1343, G1344);
nand g516(G1357, G1355, G1356);
assign G1397 = G393;
nand g518(G277, G1015, G1018);
not g519(G1019, G1015);
nand g520(G280, G1005, G1008);
not g521(G1009, G1005);
nand g522(G325, G1090, G1099);
nand g523(G364, G1189, G1192);
not g524(G1193, G1189);
nand g525(G401, G399, G400);
nand g526(G1089, G1078, G1087);
nand g527(G1139, G1137, G1138);
nand g528(G278, G1010, G1019);
nand g529(G281, G1000, G1009);
nand g530(G326, G324, G325);
nand g531(G365, G1184, G1193);
nand g532(G413, G1357, G1360);
not g533(G1361, G1357);
not g534(G1401, G1397);
nand g535(G445, G379, G918);
not g536(G1349, G1345);
nand g537(G1350, G1345, G1348);
assign G1389 = G379;
assign G1493 = G449;
assign G1501 = G449;
nand g541(G1689, G1088, G1089);
nand g542(G279, G277, G278);
nand g543(G282, G280, G281);
not g544(G1143, G1139);
nand g545(G366, G364, G365);
nand g546(G414, G1352, G1361);
nand g547(G453, G401, G918);
not g548(G1131, G1127);
nand g549(G1132, G1127, G1130);
nand g550(G1351, G1340, G1349);
not g551(G1365, G326);
assign G1405 = G401;
not g553(G285, G279);
not g554(G367, G366);
nand g555(G415, G413, G414);
not g556(G1393, G1389);
nand g557(G556, G1501, G1504);
not g558(G1505, G1501);
nand g559(G559, G1493, G1496);
not g560(G1497, G1493);
not g561(G1693, G1689);
nand g562(G1133, G1122, G1131);
assign G1477 = G445;
assign G1485 = G445;
nand g565(G1809, G1350, G1351);
not g566(G1369, G1365);
not g567(G1409, G1405);
nand g568(G557, G1498, G1505);
nand g569(G560, G1490, G1497);
assign G1362 = G282;
not g571(G1378, G415);
assign G1429 = G453;
assign G1437 = G453;
assign G1686 = G282;
nand g575(G1774, G1132, G1133);
and g576(G1910, G285, G853);
and g577(G1918, G856, G367);
nand g578(G544, G1485, G1488);
not g579(G1489, G1485);
nand g580(G547, G1477, G1480);
not g581(G1481, G1477);
nand g582(G558, G556, G557);
nand g583(G561, G559, G560);
not g584(G1813, G1809);
not g585(G1370, G348);
not g586(G1368, G1362);
not g587(G1384, G1378);
nand g588(G424, G1378, G1385);
nand g589(G508, G1437, G1440);
not g590(G1441, G1437);
nand g591(G511, G1429, G1432);
not g592(G1433, G1429);
nand g593(G545, G1482, G1489);
nand g594(G548, G1474, G1481);
not g595(G564, G558);
not g596(G1692, G1686);
nand g597(G1024, G1686, G1693);
not g598(G1780, G1774);
nand g599(G1148, G1774, G1781);
not g600(G1916, G1910);
not g601(G1924, G1918);
not g602(G1376, G1370);
nand g603(G421, G1370, G1377);
nand g604(G423, G1381, G1384);
nand g605(G509, G1434, G1441);
nand g606(G512, G1426, G1433);
nand g607(G546, G544, G545);
nand g608(G549, G547, G548);
not g609(G719, G561);
assign G722 = G561;
nand g611(G1023, G1689, G1692);
nand g612(G1147, G1777, G1780);
nand g613(G420, G1373, G1376);
nand g614(G425, G423, G424);
nand g615(G510, G508, G509);
nand g616(G513, G511, G512);
not g617(G552, G546);
nand g618(G1025, G1023, G1024);
nand g619(G1149, G1147, G1148);
not g620(G419, G418);
nand g621(G422, G420, G421);
nand g622(G441, G425, G918);
not g623(G516, G510);
not g624(G725, G549);
assign G728 = G549;
not g626(G1029, G1025);
not g627(G1153, G1149);
nand g628(G433, G419, G918);
nand g629(G437, G422, G918);
not g630(G663, G513);
assign G666 = G513;
and g632(G731, G719, G725);
and g633(G746, G722, G725);
and g634(G756, G719, G728);
and g635(G770, G722, G728);
assign G1461 = G441;
assign G1469 = G441;
assign G1413 = G433;
assign G1421 = G433;
assign G1445 = G437;
assign G1453 = G437;
nand g642(G532, G1469, G1472);
not g643(G1473, G1469);
nand g644(G535, G1461, G1464);
not g645(G1465, G1461);
nand g646(G495, G1421, G1424);
not g647(G1425, G1421);
nand g648(G498, G1413, G1416);
not g649(G1417, G1413);
not g650(G1457, G1453);
nand g651(G523, G1445, G1448);
not g652(G1449, G1445);
nand g653(G533, G1466, G1473);
nand g654(G536, G1458, G1465);
nand g655(G496, G1418, G1425);
nand g656(G499, G1410, G1417);
nand g657(G524, G1442, G1449);
nand g658(G534, G532, G533);
nand g659(G537, G535, G536);
nand g660(G497, G495, G496);
nand g661(G500, G498, G499);
nand g662(G525, G523, G524);
not g663(G540, G534);
not g664(G503, G497);
not g665(G528, G522);
not g666(G669, G537);
assign G672 = G537;
not g668(G569, G500);
and g669(G588, G566, G500);
not g670(G618, G525);
and g671(G639, G615, G525);
nand g672(G867, G516, G564, G552, G540, G482, G528, G503, G487);
assign G588a = G588;
assign G588b = G588;
assign G639a = G639;
assign G639b = G639;
and g677(G675, G663, G669);
and g678(G688, G666, G669);
and g679(G696, G663, G672);
and g680(G710, G666, G672);
and g681(G73, G949, G867, G932, G932);
and g682(G572, G565, G569);
and g683(G573, G566, G569);
and g684(G621, G614, G618);
and g685(G622, G615, G618);
nand g686(G776, G588a, G639a, G696, G731, G958);
nand g687(G780, G588a, G639a, G675, G756, G958);
nand g688(G784, G588a, G639a, G675, G746, G958);
nand g689(G788, G588a, G639a, G688, G731, G958);
nand g690(G812, G588b, G639a, G710, G746, G969);
nand g691(G832, G588b, G639b, G696, G770, G969);
nand g692(G836, G588b, G639b, G710, G756, G969);
and g693(G1509, G588a, G639a, G696, G731, G958);
and g694(G1517, G588a, G639a, G675, G756, G958);
and g695(G1525, G588a, G639a, G675, G746, G958);
and g696(G1533, G588a, G639a, G688, G731, G958);
and g697(G1581, G588b, G639a, G710, G746, G969);
and g698(G1621, G588b, G639b, G696, G770, G969);
and g699(G1629, G588b, G639b, G710, G756, G969);
nand g700(G792, G588a, G622, G696, G756, G958);
nand g701(G796, G588b, G622, G696, G746, G958);
nand g702(G800, G588b, G622, G710, G731, G958);
nand g703(G804, G588b, G622, G675, G770, G958);
nand g704(G808, G588b, G622, G688, G756, G969);
nand g705(G816, G573, G639b, G696, G756, G969);
nand g706(G820, G573, G639b, G696, G746, G969);
nand g707(G824, G573, G639b, G710, G731, G969);
nand g708(G828, G573, G639b, G688, G756, G969);
nand g709(G871, G588b, G622, G675, G731, G979);
nand g710(G873, G573, G639b, G675, G731, G979);
nand g711(G875, G573, G622, G696, G731, G979);
nand g712(G877, G573, G622, G675, G756, G979);
nand g713(G879, G573, G622, G675, G746, G979);
nand g714(G881, G573, G622, G688, G731, G979);
nand g715(G883, G573, G621, G675, G731, G979);
nand g716(G885, G572, G622, G675, G731, G979);
and g717(G1541, G588a, G622, G696, G756, G958);
and g718(G1549, G588b, G622, G696, G746, G958);
and g719(G1557, G588b, G622, G710, G731, G958);
and g720(G1565, G588b, G622, G675, G770, G958);
and g721(G1573, G588b, G622, G688, G756, G969);
and g722(G1589, G573, G639b, G696, G756, G969);
and g723(G1597, G573, G639b, G696, G746, G969);
and g724(G1605, G573, G639b, G710, G731, G969);
and g725(G1613, G573, G639b, G688, G756, G969);
nand g726(G1, G1509, G1512);
not g727(G1513, G1509);
nand g728(G4, G1517, G1520);
not g729(G1521, G1517);
nand g730(G7, G1525, G1528);
not g731(G1529, G1525);
nand g732(G10, G1533, G1536);
not g733(G1537, G1533);
nand g734(G28, G1581, G1584);
not g735(G1585, G1581);
nand g736(G43, G1621, G1624);
not g737(G1625, G1621);
nand g738(G46, G1629, G1632);
not g739(G1633, G1629);
and g740(G886, G871, G873, G875, G877, G879, G881, G883, G885);
nand g741(G2, G1506, G1513);
nand g742(G5, G1514, G1521);
nand g743(G8, G1522, G1529);
nand g744(G11, G1530, G1537);
nand g745(G13, G1541, G1544);
not g746(G1545, G1541);
nand g747(G16, G1549, G1552);
not g748(G1553, G1549);
nand g749(G19, G1557, G1560);
not g750(G1561, G1557);
nand g751(G22, G1565, G1568);
not g752(G1569, G1565);
nand g753(G25, G1573, G1576);
not g754(G1577, G1573);
nand g755(G29, G1578, G1585);
nand g756(G31, G1589, G1592);
not g757(G1593, G1589);
nand g758(G34, G1597, G1600);
not g759(G1601, G1597);
nand g760(G37, G1605, G1608);
not g761(G1609, G1605);
nand g762(G40, G1613, G1616);
not g763(G1617, G1613);
nand g764(G44, G1618, G1625);
nand g765(G47, G1626, G1633);
nand g766(G857, G776, G780, G784, G788, G792, G796, G800, G804);
nand g767(G860, G808, G812, G816, G820, G824, G828, G832, G836);
and g768(G863, G776, G780, G784, G788, G792, G796, G800, G804);
and g769(G865, G808, G812, G816, G820, G824, G828, G832, G836);
nand g770(G3, G1, G2);
nand g771(G6, G4, G5);
nand g772(G9, G7, G8);
nand g773(G12, G10, G11);
nand g774(G14, G1538, G1545);
nand g775(G17, G1546, G1553);
nand g776(G20, G1554, G1561);
nand g777(G23, G1562, G1569);
nand g778(G26, G1570, G1577);
nand g779(G30, G28, G29);
nand g780(G32, G1586, G1593);
nand g781(G35, G1594, G1601);
nand g782(G38, G1602, G1609);
nand g783(G41, G1610, G1617);
nand g784(G45, G43, G44);
nand g785(G48, G46, G47);
and g786(G1913, G857, G859);
and g787(G1921, G860, G862);
nand g788(G15, G13, G14);
nand g789(G18, G16, G17);
nand g790(G21, G19, G20);
nand g791(G24, G22, G23);
nand g792(G27, G25, G26);
nand g793(G33, G31, G32);
nand g794(G36, G34, G35);
nand g795(G39, G37, G38);
nand g796(G42, G40, G41);
and g797(G887, G863, G865, G886);
nand g798(G462, G863, G865);
and g799(G74, G949, G867, G952, G887);
nand g800(G1637, G1913, G1916);
not g801(G1917, G1913);
nand g802(G1647, G1921, G1924);
not g803(G1925, G1921);
nor g804(G75, G73, G74);
and g805(G1020, G457, G911, G462);
and g806(G1144, G469, G911, G462);
and g807(G1386, G475, G911, G462);
and g808(G1394, G478, G911, G462);
and g809(G1402, G459, G911, G462);
nand g810(G1638, G1910, G1917);
nand g811(G1648, G1918, G1925);
and g812(G1806, G472, G911, G462);
nand g813(G1639, G1637, G1638);
nand g814(G1649, G1647, G1648);
nand g815(G287, G1020, G1029);
nand g816(G350, G1144, G1153);
nand g817(G427, G1386, G1393);
nand g818(G429, G1394, G1401);
nand g819(G431, G1402, G1409);
not g820(G1028, G1020);
not g821(G1152, G1144);
not g822(G1392, G1386);
not g823(G1400, G1394);
not g824(G1408, G1402);
not g825(G1812, G1806);
nand g826(G1216, G1806, G1813);
nand g827(G286, G1025, G1028);
nand g828(G349, G1149, G1152);
nand g829(G426, G1389, G1392);
nand g830(G428, G1397, G1400);
nand g831(G430, G1405, G1408);
nand g832(G67, G1639, G1642);
not g833(G1643, G1639);
nand g834(G70, G1649, G1652);
not g835(G1653, G1649);
nand g836(G1215, G1809, G1812);
nand g837(G49, G286, G287);
nand g838(G53, G349, G350);
nand g839(G59, G426, G427);
nand g840(G61, G428, G429);
nand g841(G65, G430, G431);
nand g842(G68, G1634, G1643);
nand g843(G71, G1644, G1653);
nand g844(G1217, G1215, G1216);
and g845(G51, G49, G50);
and g846(G54, G52, G53);
and g847(G60, G58, G59);
and g848(G63, G61, G62);
and g849(G66, G64, G65);
nand g850(G69, G67, G68);
nand g851(G72, G70, G71);
nand g852(G375, G1217, G1220);
not g853(G1221, G1217);
nand g854(G376, G1212, G1221);
nand g855(G55, G375, G376);
and g856(G57, G55, G56);
not g857(in0not_0, G1362);
not g858(in1not_0, G1368);
not g859(in2not_0, G1369);
not g860(in3not_0, G1365);
and g861(T0_0, keyinput0_0, in0not_0, in1not_0, in2not_0, in3not_0);
and g862(T1_0, keyinput1_0, G1362, in1not_0, in2not_0, in3not_0);
and g863(T2_0, keyinput2_0, in0not_0, G1368, in2not_0, in3not_0);
and g864(T3_0, keyinput3_0, G1362, G1368, in2not_0, in3not_0);
and g865(T4_0, keyinput4_0, in0not_0, in1not_0, G1369, in3not_0);
and g866(T5_0, keyinput5_0, G1362, in1not_0, G1369, in3not_0);
and g867(T6_0, keyinput6_0, in0not_0, G1368, G1369, in3not_0);
and g868(T7_0, keyinput7_0, G1362, G1368, G1369, in3not_0);
and g869(T8_0, keyinput8_0, in0not_0, in1not_0, in2not_0, G1365);
and g870(T9_0, keyinput9_0, G1362, in1not_0, in2not_0, G1365);
and g871(T10_0, keyinput10_0, in0not_0, G1368, in2not_0, G1365);
and g872(T11_0, keyinput11_0, G1362, G1368, in2not_0, G1365);
and g873(T12_0, keyinput12_0, in0not_0, in1not_0, G1369, G1365);
and g874(T13_0, keyinput13_0, G1362, in1not_0, G1369, G1365);
and g875(T14_0, keyinput14_0, in0not_0, G1368, G1369, G1365);
and g876(T15_0, keyinput15_0, G1362, G1368, G1369, G1365);
or g877(G418, T0_0, T1_0, T2_0, T3_0, T4_0, T5_0, T6_0, T7_0, T8_0, T9_0, T10_0, T11_0, T12_0, T13_0, T14_0, T15_0);
not g878(in0not_1, G989);
not g879(in1not_1, G985);
not g880(in2not_1, G988);
not g881(in3not_1, G980);
and g882(T0_1, keyinput0_1, in0not_1, in1not_1, in2not_1, in3not_1);
and g883(T1_1, keyinput1_1, G989, in1not_1, in2not_1, in3not_1);
and g884(T2_1, keyinput2_1, in0not_1, G985, in2not_1, in3not_1);
and g885(T3_1, keyinput3_1, G989, G985, in2not_1, in3not_1);
and g886(T4_1, keyinput4_1, in0not_1, in1not_1, G988, in3not_1);
and g887(T5_1, keyinput5_1, G989, in1not_1, G988, in3not_1);
and g888(T6_1, keyinput6_1, in0not_1, G985, G988, in3not_1);
and g889(T7_1, keyinput7_1, G989, G985, G988, in3not_1);
and g890(T8_1, keyinput8_1, in0not_1, in1not_1, in2not_1, G980);
and g891(T9_1, keyinput9_1, G989, in1not_1, in2not_1, G980);
and g892(T10_1, keyinput10_1, in0not_1, G985, in2not_1, G980);
and g893(T11_1, keyinput11_1, G989, G985, in2not_1, G980);
and g894(T12_1, keyinput12_1, in0not_1, in1not_1, G988, G980);
and g895(T13_1, keyinput13_1, G989, in1not_1, G988, G980);
and g896(T14_1, keyinput14_1, in0not_1, G985, G988, G980);
and g897(T15_1, keyinput15_1, G989, G985, G988, G980);
or g898(G262, T0_1, T1_1, T2_1, T3_1, T4_1, T5_1, T6_1, T7_1, T8_1, T9_1, T10_1, T11_1, T12_1, T13_1, T14_1, T15_1);
not g899(in0not_2, G1139);
not g900(in1not_2, G1142);
not g901(in2not_2, G1143);
not g902(in3not_2, G1134);
and g903(T0_2, keyinput0_2, in0not_2, in1not_2, in2not_2, in3not_2);
and g904(T1_2, keyinput1_2, G1139, in1not_2, in2not_2, in3not_2);
and g905(T2_2, keyinput2_2, in0not_2, G1142, in2not_2, in3not_2);
and g906(T3_2, keyinput3_2, G1139, G1142, in2not_2, in3not_2);
and g907(T4_2, keyinput4_2, in0not_2, in1not_2, G1143, in3not_2);
and g908(T5_2, keyinput5_2, G1139, in1not_2, G1143, in3not_2);
and g909(T6_2, keyinput6_2, in0not_2, G1142, G1143, in3not_2);
and g910(T7_2, keyinput7_2, G1139, G1142, G1143, in3not_2);
and g911(T8_2, keyinput8_2, in0not_2, in1not_2, in2not_2, G1134);
and g912(T9_2, keyinput9_2, G1139, in1not_2, in2not_2, G1134);
and g913(T10_2, keyinput10_2, in0not_2, G1142, in2not_2, G1134);
and g914(T11_2, keyinput11_2, G1139, G1142, in2not_2, G1134);
and g915(T12_2, keyinput12_2, in0not_2, in1not_2, G1143, G1134);
and g916(T13_2, keyinput13_2, G1139, in1not_2, G1143, G1134);
and g917(T14_2, keyinput14_2, in0not_2, G1142, G1143, G1134);
and g918(T15_2, keyinput15_2, G1139, G1142, G1143, G1134);
or g919(G348, T0_2, T1_2, T2_2, T3_2, T4_2, T5_2, T6_2, T7_2, T8_2, T9_2, T10_2, T11_2, T12_2, T13_2, T14_2, T15_2);
not g920(in0not_3, G1765);
not g921(in1not_3, G1764);
not g922(in2not_3, G1758);
not g923(in3not_3, G1761);
and g924(T0_3, keyinput0_3, in0not_3, in1not_3, in2not_3, in3not_3);
and g925(T1_3, keyinput1_3, G1765, in1not_3, in2not_3, in3not_3);
and g926(T2_3, keyinput2_3, in0not_3, G1764, in2not_3, in3not_3);
and g927(T3_3, keyinput3_3, G1765, G1764, in2not_3, in3not_3);
and g928(T4_3, keyinput4_3, in0not_3, in1not_3, G1758, in3not_3);
and g929(T5_3, keyinput5_3, G1765, in1not_3, G1758, in3not_3);
and g930(T6_3, keyinput6_3, in0not_3, G1764, G1758, in3not_3);
and g931(T7_3, keyinput7_3, G1765, G1764, G1758, in3not_3);
and g932(T8_3, keyinput8_3, in0not_3, in1not_3, in2not_3, G1761);
and g933(T9_3, keyinput9_3, G1765, in1not_3, in2not_3, G1761);
and g934(T10_3, keyinput10_3, in0not_3, G1764, in2not_3, G1761);
and g935(T11_3, keyinput11_3, G1765, G1764, in2not_3, G1761);
and g936(T12_3, keyinput12_3, in0not_3, in1not_3, G1758, G1761);
and g937(T13_3, keyinput13_3, G1765, in1not_3, G1758, G1761);
and g938(T14_3, keyinput14_3, in0not_3, G1764, G1758, G1761);
and g939(T15_3, keyinput15_3, G1765, G1764, G1758, G1761);
or g940(G1127, T0_3, T1_3, T2_3, T3_3, T4_3, T5_3, T6_3, T7_3, T8_3, T9_3, T10_3, T11_3, T12_3, T13_3, T14_3, T15_3);
not g941(in0not_4, G1457);
not g942(in1not_4, G1453);
not g943(in2not_4, G1456);
not g944(in3not_4, G1450);
and g945(T0_4, keyinput0_4, in0not_4, in1not_4, in2not_4, in3not_4);
and g946(T1_4, keyinput1_4, G1457, in1not_4, in2not_4, in3not_4);
and g947(T2_4, keyinput2_4, in0not_4, G1453, in2not_4, in3not_4);
and g948(T3_4, keyinput3_4, G1457, G1453, in2not_4, in3not_4);
and g949(T4_4, keyinput4_4, in0not_4, in1not_4, G1456, in3not_4);
and g950(T5_4, keyinput5_4, G1457, in1not_4, G1456, in3not_4);
and g951(T6_4, keyinput6_4, in0not_4, G1453, G1456, in3not_4);
and g952(T7_4, keyinput7_4, G1457, G1453, G1456, in3not_4);
and g953(T8_4, keyinput8_4, in0not_4, in1not_4, in2not_4, G1450);
and g954(T9_4, keyinput9_4, G1457, in1not_4, in2not_4, G1450);
and g955(T10_4, keyinput10_4, in0not_4, G1453, in2not_4, G1450);
and g956(T11_4, keyinput11_4, G1457, G1453, in2not_4, G1450);
and g957(T12_4, keyinput12_4, in0not_4, in1not_4, G1456, G1450);
and g958(T13_4, keyinput13_4, G1457, in1not_4, G1456, G1450);
and g959(T14_4, keyinput14_4, in0not_4, G1453, G1456, G1450);
and g960(T15_4, keyinput15_4, G1457, G1453, G1456, G1450);
or g961(G522, T0_4, T1_4, T2_4, T3_4, T4_4, T5_4, T6_4, T7_4, T8_4, T9_4, T10_4, T11_4, T12_4, T13_4, T14_4, T15_4);
not g962(in0not_5, G1885);
not g963(in1not_5, G1884);
not g964(in2not_5, G1881);
not g965(in3not_5, G1878);
and g966(T0_5, keyinput0_5, in0not_5, in1not_5, in2not_5, in3not_5);
and g967(T1_5, keyinput1_5, G1885, in1not_5, in2not_5, in3not_5);
and g968(T2_5, keyinput2_5, in0not_5, G1884, in2not_5, in3not_5);
and g969(T3_5, keyinput3_5, G1885, G1884, in2not_5, in3not_5);
and g970(T4_5, keyinput4_5, in0not_5, in1not_5, G1881, in3not_5);
and g971(T5_5, keyinput5_5, G1885, in1not_5, G1881, in3not_5);
and g972(T6_5, keyinput6_5, in0not_5, G1884, G1881, in3not_5);
and g973(T7_5, keyinput7_5, G1885, G1884, G1881, in3not_5);
and g974(T8_5, keyinput8_5, in0not_5, in1not_5, in2not_5, G1878);
and g975(T9_5, keyinput9_5, G1885, in1not_5, in2not_5, G1878);
and g976(T10_5, keyinput10_5, in0not_5, G1884, in2not_5, G1878);
and g977(T11_5, keyinput11_5, G1885, G1884, in2not_5, G1878);
and g978(T12_5, keyinput12_5, in0not_5, in1not_5, G1881, G1878);
and g979(T13_5, keyinput13_5, G1885, in1not_5, G1881, G1878);
and g980(T14_5, keyinput14_5, in0not_5, G1884, G1881, G1878);
and g981(T15_5, keyinput15_5, G1885, G1884, G1881, G1878);
or g982(G1317, T0_5, T1_5, T2_5, T3_5, T4_5, T5_5, T6_5, T7_5, T8_5, T9_5, T10_5, T11_5, T12_5, T13_5, T14_5, T15_5);
not g983(in0not_6, G943);
not g984(in1not_6, G893);
not g985(in2not_6, G919);
not g986(in3not_6, G907);
and g987(T0_6, keyinput0_6, in0not_6, in1not_6, in2not_6, in3not_6);
and g988(T1_6, keyinput1_6, G943, in1not_6, in2not_6, in3not_6);
and g989(T2_6, keyinput2_6, in0not_6, G893, in2not_6, in3not_6);
and g990(T3_6, keyinput3_6, G943, G893, in2not_6, in3not_6);
and g991(T4_6, keyinput4_6, in0not_6, in1not_6, G919, in3not_6);
and g992(T5_6, keyinput5_6, G943, in1not_6, G919, in3not_6);
and g993(T6_6, keyinput6_6, in0not_6, G893, G919, in3not_6);
and g994(T7_6, keyinput7_6, G943, G893, G919, in3not_6);
and g995(T8_6, keyinput8_6, in0not_6, in1not_6, in2not_6, G907);
and g996(T9_6, keyinput9_6, G943, in1not_6, in2not_6, G907);
and g997(T10_6, keyinput10_6, in0not_6, G893, in2not_6, G907);
and g998(T11_6, keyinput11_6, G943, G893, in2not_6, G907);
and g999(T12_6, keyinput12_6, in0not_6, in1not_6, G919, G907);
and g1000(T13_6, keyinput13_6, G943, in1not_6, G919, G907);
and g1001(T14_6, keyinput14_6, in0not_6, G893, G919, G907);
and g1002(T15_6, keyinput15_6, G943, G893, G919, G907);
or g1003(G956, T0_6, T1_6, T2_6, T3_6, T4_6, T5_6, T6_6, T7_6, T8_6, T9_6, T10_6, T11_6, T12_6, T13_6, T14_6, T15_6);
not g1004(in0not_7, G1121);
not g1005(in1not_7, G1117);
not g1006(in2not_7, G1120);
not g1007(in3not_7, G1112);
and g1008(T0_7, keyinput0_7, in0not_7, in1not_7, in2not_7, in3not_7);
and g1009(T1_7, keyinput1_7, G1121, in1not_7, in2not_7, in3not_7);
and g1010(T2_7, keyinput2_7, in0not_7, G1117, in2not_7, in3not_7);
and g1011(T3_7, keyinput3_7, G1121, G1117, in2not_7, in3not_7);
and g1012(T4_7, keyinput4_7, in0not_7, in1not_7, G1120, in3not_7);
and g1013(T5_7, keyinput5_7, G1121, in1not_7, G1120, in3not_7);
and g1014(T6_7, keyinput6_7, in0not_7, G1117, G1120, in3not_7);
and g1015(T7_7, keyinput7_7, G1121, G1117, G1120, in3not_7);
and g1016(T8_7, keyinput8_7, in0not_7, in1not_7, in2not_7, G1112);
and g1017(T9_7, keyinput9_7, G1121, in1not_7, in2not_7, G1112);
and g1018(T10_7, keyinput10_7, in0not_7, G1117, in2not_7, G1112);
and g1019(T11_7, keyinput11_7, G1121, G1117, in2not_7, G1112);
and g1020(T12_7, keyinput12_7, in0not_7, in1not_7, G1120, G1112);
and g1021(T13_7, keyinput13_7, G1121, in1not_7, G1120, G1112);
and g1022(T14_7, keyinput14_7, in0not_7, G1117, G1120, G1112);
and g1023(T15_7, keyinput15_7, G1121, G1117, G1120, G1112);
or g1024(G336, T0_7, T1_7, T2_7, T3_7, T4_7, T5_7, T6_7, T7_7, T8_7, T9_7, T10_7, T11_7, T12_7, T13_7, T14_7, T15_7);
endmodule
