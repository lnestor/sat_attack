
module c3540 ( N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, 
        N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, 
        N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, 
        N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, 
        N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, 
        N4815, N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, 
        N5231, N5360, N5361, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116,
         N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190,
         N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264,
         N270, N274, N283, N294, N303, N311, N317, N322, N326, N329, N330,
         N343, N349, N350, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815,
         N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231,
         N5360, N5361;
  wire   n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286;

  NAND2X0 U654 ( .IN1(n640), .IN2(n641), .QN(N5361) );
  XOR2X1 U655 ( .IN1(keyinput127), .IN2(n642), .Q(n641) );
  NOR2X0 U656 ( .IN1(n643), .IN2(n644), .QN(n642) );
  XOR2X1 U657 ( .IN1(keyinput125), .IN2(n645), .Q(n644) );
  XOR2X1 U658 ( .IN1(n646), .IN2(n647), .Q(n643) );
  XOR2X1 U659 ( .IN1(n648), .IN2(n645), .Q(n640) );
  XNOR2X1 U660 ( .IN1(n649), .IN2(n650), .Q(n645) );
  NOR2X0 U661 ( .IN1(n651), .IN2(n652), .QN(n650) );
  XOR2X1 U662 ( .IN1(keyinput119), .IN2(n653), .Q(n652) );
  NAND2X0 U663 ( .IN1(n654), .IN2(keyinput126), .QN(n648) );
  XOR2X1 U664 ( .IN1(n655), .IN2(n647), .Q(n654) );
  MUX21X1 U665 ( .IN1(n656), .IN2(n657), .S(n658), .Q(N5360) );
  OA21X1 U666 ( .IN1(n646), .IN2(n659), .IN3(n660), .Q(n658) );
  MUX21X1 U667 ( .IN1(n661), .IN2(n662), .S(n647), .Q(n660) );
  OA21X1 U668 ( .IN1(n663), .IN2(N5078), .IN3(n664), .Q(n647) );
  XNOR2X1 U669 ( .IN1(n665), .IN2(keyinput118), .Q(n664) );
  NAND2X0 U670 ( .IN1(N5078), .IN2(n663), .QN(n665) );
  NAND2X0 U671 ( .IN1(n646), .IN2(n659), .QN(n662) );
  NOR2X0 U672 ( .IN1(keyinput122), .IN2(n666), .QN(n661) );
  XOR2X1 U673 ( .IN1(keyinput121), .IN2(n646), .Q(n666) );
  INVX0 U674 ( .INP(keyinput122), .ZN(n659) );
  INVX0 U675 ( .INP(n655), .ZN(n646) );
  NAND2X0 U676 ( .IN1(n667), .IN2(n668), .QN(n655) );
  AO21X1 U677 ( .IN1(keyinput117), .IN2(N4815), .IN3(N5047), .Q(n668) );
  MUX21X1 U678 ( .IN1(keyinput114), .IN2(n669), .S(N4815), .Q(n667) );
  NAND3X0 U679 ( .IN1(keyinput114), .IN2(N5047), .IN3(keyinput117), .QN(n669)
         );
  AO21X1 U680 ( .IN1(keyinput123), .IN2(n670), .IN3(n671), .Q(n657) );
  NOR3X0 U681 ( .IN1(n670), .IN2(keyinput123), .IN3(n671), .QN(n656) );
  MUX21X1 U682 ( .IN1(n649), .IN2(n672), .S(n673), .Q(n671) );
  XNOR2X1 U683 ( .IN1(n674), .IN2(n675), .Q(n673) );
  OA21X1 U684 ( .IN1(n651), .IN2(n653), .IN3(n676), .Q(n675) );
  XOR2X1 U685 ( .IN1(keyinput16), .IN2(n677), .Q(n676) );
  NOR2X0 U686 ( .IN1(n678), .IN2(N5102), .QN(n653) );
  NOR2X0 U687 ( .IN1(n679), .IN2(N5120), .QN(n651) );
  NAND2X0 U688 ( .IN1(N350), .IN2(n677), .QN(n674) );
  AND2X1 U689 ( .IN1(N213), .IN2(n680), .Q(n677) );
  AOI21X1 U690 ( .IN1(N5121), .IN2(N4944), .IN3(n681), .QN(n672) );
  NAND2X0 U691 ( .IN1(n682), .IN2(n683), .QN(n649) );
  INVX0 U692 ( .INP(n681), .ZN(n683) );
  MUX21X1 U693 ( .IN1(n684), .IN2(N5121), .S(keyinput120), .Q(n682) );
  NAND2X0 U694 ( .IN1(N4944), .IN2(N5121), .QN(n684) );
  INVX0 U695 ( .INP(keyinput124), .ZN(n670) );
  NAND3X0 U696 ( .IN1(n685), .IN2(N5192), .IN3(N213), .QN(N5231) );
  NAND3X0 U697 ( .IN1(n678), .IN2(n680), .IN3(n679), .QN(n685) );
  INVX0 U698 ( .INP(N5102), .ZN(n679) );
  INVX0 U699 ( .INP(N343), .ZN(n680) );
  INVX0 U700 ( .INP(N5120), .ZN(n678) );
  NAND4X0 U701 ( .IN1(n686), .IN2(n663), .IN3(n681), .IN4(n687), .QN(N5192) );
  NOR4X0 U702 ( .IN1(N5120), .IN2(N5078), .IN3(N5102), .IN4(N5047), .QN(n687)
         );
  NOR2X0 U703 ( .IN1(N4944), .IN2(N5121), .QN(n681) );
  INVX0 U704 ( .INP(N5045), .ZN(n663) );
  AO222X1 U705 ( .IN1(n688), .IN2(n689), .IN3(n690), .IN4(n691), .IN5(n692), 
        .IN6(n693), .Q(N5121) );
  OA221X1 U706 ( .IN1(n694), .IN2(n695), .IN3(N68), .IN4(n696), .IN5(n697), 
        .Q(n691) );
  NAND4X0 U707 ( .IN1(n698), .IN2(n699), .IN3(n700), .IN4(n701), .QN(n697) );
  OA221X1 U708 ( .IN1(n702), .IN2(n703), .IN3(n704), .IN4(n705), .IN5(n706), 
        .Q(n701) );
  OA222X1 U709 ( .IN1(n707), .IN2(n708), .IN3(n709), .IN4(n710), .IN5(n711), 
        .IN6(n712), .Q(n706) );
  XNOR2X1 U710 ( .IN1(keyinput55), .IN2(n713), .Q(n710) );
  OA22X1 U711 ( .IN1(n714), .IN2(n715), .IN3(n716), .IN4(n717), .Q(n700) );
  XOR2X1 U712 ( .IN1(n718), .IN2(keyinput68), .Q(n698) );
  NAND2X0 U713 ( .IN1(n719), .IN2(N159), .QN(n718) );
  XNOR2X1 U714 ( .IN1(n720), .IN2(keyinput80), .Q(n695) );
  NAND4X0 U715 ( .IN1(n721), .IN2(N33), .IN3(n722), .IN4(n723), .QN(n720) );
  OA221X1 U716 ( .IN1(n724), .IN2(n703), .IN3(n713), .IN4(n725), .IN5(n726), 
        .Q(n723) );
  OA222X1 U717 ( .IN1(n704), .IN2(n727), .IN3(n711), .IN4(n728), .IN5(n707), 
        .IN6(n729), .Q(n726) );
  OA22X1 U718 ( .IN1(n714), .IN2(n730), .IN3(n731), .IN4(n732), .Q(n722) );
  XOR2X1 U719 ( .IN1(n733), .IN2(keyinput72), .Q(n721) );
  NAND2X0 U720 ( .IN1(N87), .IN2(n734), .QN(n733) );
  NOR2X0 U721 ( .IN1(n735), .IN2(n736), .QN(n690) );
  XOR2X1 U722 ( .IN1(n737), .IN2(keyinput98), .Q(n735) );
  NAND2X0 U723 ( .IN1(n738), .IN2(n739), .QN(n737) );
  XOR2X1 U724 ( .IN1(n692), .IN2(n740), .Q(n688) );
  AO221X1 U725 ( .IN1(n741), .IN2(n689), .IN3(n742), .IN4(n693), .IN5(n743), 
        .Q(N5120) );
  OA221X1 U726 ( .IN1(N50), .IN2(n696), .IN3(n694), .IN4(n744), .IN5(n745), 
        .Q(n743) );
  OA21X1 U727 ( .IN1(n746), .IN2(n747), .IN3(n748), .Q(n745) );
  MUX21X1 U728 ( .IN1(n749), .IN2(N50), .S(N41), .Q(n744) );
  MUX21X1 U729 ( .IN1(n750), .IN2(n751), .S(N33), .Q(n749) );
  NAND4X0 U730 ( .IN1(n752), .IN2(n753), .IN3(n754), .IN4(n755), .QN(n751) );
  OA22X1 U731 ( .IN1(n756), .IN2(n757), .IN3(n731), .IN4(n711), .Q(n755) );
  XOR2X1 U732 ( .IN1(n716), .IN2(keyinput59), .Q(n756) );
  OA22X1 U733 ( .IN1(n707), .IN2(n758), .IN3(n704), .IN4(n729), .Q(n754) );
  OA22X1 U734 ( .IN1(n713), .IN2(n728), .IN3(n702), .IN4(n703), .Q(n753) );
  OA22X1 U735 ( .IN1(n714), .IN2(n727), .IN3(n724), .IN4(n732), .Q(n752) );
  NAND4X0 U736 ( .IN1(n759), .IN2(n760), .IN3(n761), .IN4(n762), .QN(n750) );
  AOI22X1 U737 ( .IN1(N124), .IN2(n763), .IN3(N143), .IN4(n764), .QN(n762) );
  XOR2X1 U738 ( .IN1(keyinput52), .IN2(n719), .Q(n764) );
  XOR2X1 U739 ( .IN1(keyinput51), .IN2(n765), .Q(n763) );
  OA22X1 U740 ( .IN1(n711), .IN2(n709), .IN3(n707), .IN4(n705), .Q(n761) );
  OA22X1 U741 ( .IN1(n704), .IN2(n715), .IN3(n713), .IN4(n766), .Q(n760) );
  OA22X1 U742 ( .IN1(n703), .IN2(n767), .IN3(n716), .IN4(n708), .Q(n759) );
  MUX21X1 U743 ( .IN1(n768), .IN2(n769), .S(n740), .Q(n741) );
  AND3X1 U744 ( .IN1(n770), .IN2(n692), .IN3(n742), .Q(n769) );
  XOR2X1 U745 ( .IN1(n771), .IN2(n772), .Q(n742) );
  NAND2X0 U746 ( .IN1(keyinput112), .IN2(n773), .QN(n771) );
  AO21X1 U747 ( .IN1(n773), .IN2(n772), .IN3(n774), .Q(n768) );
  XOR2X1 U748 ( .IN1(n775), .IN2(keyinput115), .Q(n774) );
  OR2X1 U749 ( .IN1(n772), .IN2(n773), .Q(n775) );
  XNOR2X1 U750 ( .IN1(n776), .IN2(n777), .Q(n773) );
  NAND2X0 U751 ( .IN1(keyinput110), .IN2(n747), .QN(n776) );
  XOR2X1 U752 ( .IN1(n778), .IN2(n779), .Q(n747) );
  NAND2X0 U753 ( .IN1(n780), .IN2(n781), .QN(n778) );
  AO221X1 U754 ( .IN1(n689), .IN2(n782), .IN3(n783), .IN4(n693), .IN5(n784), 
        .Q(N5078) );
  XNOR2X1 U755 ( .IN1(n785), .IN2(keyinput103), .Q(n784) );
  NAND4X0 U756 ( .IN1(n748), .IN2(n786), .IN3(n787), .IN4(n788), .QN(n785) );
  NAND4X0 U757 ( .IN1(n699), .IN2(n789), .IN3(n790), .IN4(n791), .QN(n788) );
  OA221X1 U758 ( .IN1(n757), .IN2(n732), .IN3(n716), .IN4(n724), .IN5(n792), 
        .Q(n791) );
  OA222X1 U759 ( .IN1(n714), .IN2(n712), .IN3(n707), .IN4(n702), .IN5(n703), 
        .IN6(n758), .Q(n792) );
  OA22X1 U760 ( .IN1(n711), .IN2(n717), .IN3(n704), .IN4(n767), .Q(n790) );
  OR2X1 U761 ( .IN1(n708), .IN2(n713), .Q(n789) );
  OA21X1 U762 ( .IN1(n793), .IN2(n794), .IN3(n795), .Q(n787) );
  NAND3X0 U763 ( .IN1(n796), .IN2(n797), .IN3(n798), .QN(n795) );
  XNOR2X1 U764 ( .IN1(keyinput96), .IN2(n799), .Q(n796) );
  OA221X1 U765 ( .IN1(N97), .IN2(n800), .IN3(n801), .IN4(n802), .IN5(n803), 
        .Q(n793) );
  XOR2X1 U766 ( .IN1(keyinput33), .IN2(n804), .Q(n802) );
  NAND4X0 U767 ( .IN1(n805), .IN2(n806), .IN3(n807), .IN4(n808), .QN(n786) );
  OA221X1 U768 ( .IN1(n732), .IN2(n727), .IN3(n714), .IN4(n809), .IN5(n810), 
        .Q(n808) );
  OA222X1 U769 ( .IN1(n703), .IN2(n729), .IN3(n707), .IN4(n725), .IN5(n704), 
        .IN6(n811), .Q(n810) );
  OA21X1 U770 ( .IN1(n713), .IN2(n812), .IN3(n813), .Q(n807) );
  XOR2X1 U771 ( .IN1(n814), .IN2(keyinput73), .Q(n806) );
  NAND2X0 U772 ( .IN1(N116), .IN2(n734), .QN(n814) );
  XOR2X1 U773 ( .IN1(n815), .IN2(keyinput74), .Q(n805) );
  NAND2X0 U774 ( .IN1(N303), .IN2(n816), .QN(n815) );
  INVX0 U775 ( .INP(n817), .ZN(n783) );
  XOR2X1 U776 ( .IN1(n818), .IN2(n817), .Q(n782) );
  NAND2X0 U777 ( .IN1(n819), .IN2(n820), .QN(n818) );
  NAND2X0 U778 ( .IN1(n821), .IN2(n822), .QN(N5102) );
  NAND3X0 U779 ( .IN1(n748), .IN2(n823), .IN3(n824), .QN(n822) );
  AOI222X1 U780 ( .IN1(n825), .IN2(n826), .IN3(n827), .IN4(n828), .IN5(n829), 
        .IN6(n830), .QN(n824) );
  OA221X1 U781 ( .IN1(n757), .IN2(n703), .IN3(n713), .IN4(n727), .IN5(n831), 
        .Q(n828) );
  OA222X1 U782 ( .IN1(n731), .IN2(n707), .IN3(n832), .IN4(n728), .IN5(n711), 
        .IN6(n729), .Q(n831) );
  XOR2X1 U783 ( .IN1(n833), .IN2(keyinput60), .Q(n832) );
  OA221X1 U784 ( .IN1(n716), .IN2(n724), .IN3(n714), .IN4(n725), .IN5(n834), 
        .Q(n827) );
  OA21X1 U785 ( .IN1(n732), .IN2(n758), .IN3(n813), .Q(n834) );
  OA221X1 U786 ( .IN1(n704), .IN2(n709), .IN3(n707), .IN4(n712), .IN5(n835), 
        .Q(n826) );
  OA222X1 U787 ( .IN1(n711), .IN2(n705), .IN3(n766), .IN4(n836), .IN5(n715), 
        .IN6(n837), .Q(n835) );
  XNOR2X1 U788 ( .IN1(keyinput54), .IN2(n713), .Q(n837) );
  INVX0 U789 ( .INP(N128), .ZN(n715) );
  XOR2X1 U790 ( .IN1(keyinput53), .IN2(n765), .Q(n836) );
  INVX0 U791 ( .INP(N125), .ZN(n766) );
  OA221X1 U792 ( .IN1(n716), .IN2(n767), .IN3(n717), .IN4(n703), .IN5(n838), 
        .Q(n825) );
  OA21X1 U793 ( .IN1(n732), .IN2(n708), .IN3(n699), .Q(n838) );
  NAND2X0 U794 ( .IN1(n839), .IN2(n739), .QN(n823) );
  XOR2X1 U795 ( .IN1(n840), .IN2(n841), .Q(n839) );
  MUX21X1 U796 ( .IN1(n842), .IN2(n843), .S(n770), .Q(n821) );
  XOR3X1 U797 ( .IN1(n844), .IN2(n845), .IN3(n846), .Q(n770) );
  NOR2X0 U798 ( .IN1(n847), .IN2(keyinput104), .QN(n844) );
  OA22X1 U799 ( .IN1(n848), .IN2(n738), .IN3(n849), .IN4(n850), .Q(n847) );
  OA21X1 U800 ( .IN1(n851), .IN2(n852), .IN3(n853), .Q(n843) );
  XOR2X1 U801 ( .IN1(n693), .IN2(keyinput32), .Q(n853) );
  NOR2X0 U802 ( .IN1(n854), .IN2(n855), .QN(n851) );
  OR3X1 U803 ( .IN1(n852), .IN2(n854), .IN3(n855), .Q(n842) );
  INVX0 U804 ( .INP(n740), .ZN(n855) );
  NOR2X0 U805 ( .IN1(n856), .IN2(n857), .QN(n740) );
  NOR3X0 U806 ( .IN1(keyinput108), .IN2(n858), .IN3(n859), .QN(n857) );
  INVX0 U807 ( .INP(n692), .ZN(n854) );
  AO21X1 U808 ( .IN1(n846), .IN2(n860), .IN3(n861), .Q(n692) );
  MUX21X1 U809 ( .IN1(n862), .IN2(n863), .S(n864), .Q(n861) );
  NOR2X0 U810 ( .IN1(n865), .IN2(n860), .QN(n863) );
  XOR2X1 U811 ( .IN1(n860), .IN2(n865), .Q(n862) );
  INVX0 U812 ( .INP(n848), .ZN(n860) );
  OA22X1 U813 ( .IN1(n866), .IN2(n849), .IN3(n867), .IN4(n868), .Q(n848) );
  XNOR2X1 U814 ( .IN1(n869), .IN2(keyinput49), .Q(n852) );
  AO222X1 U815 ( .IN1(n689), .IN2(n870), .IN3(n871), .IN4(n872), .IN5(n820), 
        .IN6(n693), .Q(N5047) );
  OA221X1 U816 ( .IN1(n873), .IN2(n874), .IN3(n875), .IN4(n876), .IN5(n877), 
        .Q(n872) );
  NAND4X0 U817 ( .IN1(n878), .IN2(n699), .IN3(n879), .IN4(n880), .QN(n877) );
  OA221X1 U818 ( .IN1(n714), .IN2(n708), .IN3(n731), .IN4(n703), .IN5(n881), 
        .Q(n880) );
  OA222X1 U819 ( .IN1(n713), .IN2(n767), .IN3(n882), .IN4(n702), .IN5(n704), 
        .IN6(n717), .Q(n881) );
  XOR2X1 U820 ( .IN1(n711), .IN2(keyinput58), .Q(n882) );
  OA22X1 U821 ( .IN1(n716), .IN2(n758), .IN3(n724), .IN4(n732), .Q(n879) );
  XOR2X1 U822 ( .IN1(n883), .IN2(keyinput71), .Q(n878) );
  NAND2X0 U823 ( .IN1(n884), .IN2(N68), .QN(n883) );
  XNOR2X1 U824 ( .IN1(n885), .IN2(keyinput76), .Q(n874) );
  NAND4X0 U825 ( .IN1(n886), .IN2(n887), .IN3(n888), .IN4(n889), .QN(n885) );
  OA221X1 U826 ( .IN1(n711), .IN2(n811), .IN3(n890), .IN4(n725), .IN5(n891), 
        .Q(n889) );
  OA22X1 U827 ( .IN1(n707), .IN2(n730), .IN3(n704), .IN4(n812), .Q(n891) );
  XOR2X1 U828 ( .IN1(n732), .IN2(keyinput64), .Q(n890) );
  OA22X1 U829 ( .IN1(n713), .IN2(n809), .IN3(n714), .IN4(n892), .Q(n888) );
  NAND2X0 U830 ( .IN1(N283), .IN2(n734), .QN(n887) );
  XOR2X1 U831 ( .IN1(keyinput75), .IN2(n893), .Q(n886) );
  NOR2X0 U832 ( .IN1(n703), .IN2(n728), .QN(n893) );
  OA21X1 U833 ( .IN1(n894), .IN2(n794), .IN3(n748), .Q(n871) );
  OA221X1 U834 ( .IN1(N107), .IN2(n895), .IN3(n896), .IN4(n803), .IN5(n897), 
        .Q(n894) );
  XOR2X1 U835 ( .IN1(n898), .IN2(keyinput85), .Q(n897) );
  NAND2X0 U836 ( .IN1(n899), .IN2(n900), .QN(n898) );
  XOR2X1 U837 ( .IN1(n901), .IN2(keyinput34), .Q(n900) );
  MUX21X1 U838 ( .IN1(n902), .IN2(n903), .S(n904), .Q(n899) );
  NAND4X0 U839 ( .IN1(n896), .IN2(N58), .IN3(n905), .IN4(n717), .QN(n903) );
  NAND2X0 U840 ( .IN1(N77), .IN2(N68), .QN(n905) );
  XOR2X1 U841 ( .IN1(n906), .IN2(n907), .Q(n902) );
  INVX0 U842 ( .INP(n908), .ZN(n896) );
  XOR2X1 U843 ( .IN1(keyinput35), .IN2(n909), .Q(n895) );
  XOR3X1 U844 ( .IN1(n819), .IN2(n910), .IN3(n911), .Q(n870) );
  NAND2X0 U845 ( .IN1(keyinput102), .IN2(n912), .QN(n911) );
  AO221X1 U846 ( .IN1(n913), .IN2(n914), .IN3(n915), .IN4(n693), .IN5(n916), 
        .Q(N5045) );
  XOR2X1 U847 ( .IN1(keyinput116), .IN2(n917), .Q(n916) );
  NOR2X0 U848 ( .IN1(n918), .IN2(n869), .QN(n917) );
  OA22X1 U849 ( .IN1(n817), .IN2(n919), .IN3(n819), .IN4(n920), .Q(n918) );
  XOR2X1 U850 ( .IN1(n921), .IN2(n922), .Q(n920) );
  INVX0 U851 ( .INP(n923), .ZN(n819) );
  AO21X1 U852 ( .IN1(n924), .IN2(n925), .IN3(n926), .Q(n919) );
  INVX0 U853 ( .INP(n820), .ZN(n926) );
  AO21X1 U854 ( .IN1(n912), .IN2(n910), .IN3(n927), .Q(n820) );
  XOR2X1 U855 ( .IN1(keyinput111), .IN2(n928), .Q(n927) );
  NOR2X0 U856 ( .IN1(n912), .IN2(n910), .QN(n928) );
  XOR2X1 U857 ( .IN1(n875), .IN2(n929), .Q(n912) );
  OR3X1 U858 ( .IN1(n923), .IN2(keyinput113), .IN3(n921), .Q(n925) );
  XOR2X1 U859 ( .IN1(n930), .IN2(n931), .Q(n817) );
  OA21X1 U860 ( .IN1(n932), .IN2(n933), .IN3(keyinput107), .Q(n931) );
  XOR2X1 U861 ( .IN1(n934), .IN2(keyinput109), .Q(n933) );
  NAND2X0 U862 ( .IN1(n935), .IN2(n936), .QN(n934) );
  NOR2X0 U863 ( .IN1(n935), .IN2(n936), .QN(n932) );
  OAI21X1 U864 ( .IN1(n921), .IN2(keyinput113), .IN3(n924), .QN(n915) );
  MUX21X1 U865 ( .IN1(n922), .IN2(n937), .S(n921), .Q(n924) );
  NAND2X0 U866 ( .IN1(keyinput113), .IN2(n922), .QN(n937) );
  INVX0 U867 ( .INP(n938), .ZN(n922) );
  MUX21X1 U868 ( .IN1(n939), .IN2(n940), .S(keyinput100), .Q(n938) );
  OR2X1 U869 ( .IN1(n930), .IN2(n941), .Q(n940) );
  NAND2X0 U870 ( .IN1(N330), .IN2(n942), .QN(n939) );
  NAND3X0 U871 ( .IN1(n943), .IN2(n936), .IN3(n875), .QN(n942) );
  AO21X1 U872 ( .IN1(n944), .IN2(n945), .IN3(n946), .Q(n921) );
  MUX21X1 U873 ( .IN1(n947), .IN2(n948), .S(n949), .Q(n946) );
  NOR2X0 U874 ( .IN1(n947), .IN2(n945), .QN(n948) );
  NAND2X0 U875 ( .IN1(keyinput99), .IN2(n950), .QN(n947) );
  INVX0 U876 ( .INP(n944), .ZN(n950) );
  INVX0 U877 ( .INP(keyinput106), .ZN(n945) );
  OA22X1 U878 ( .IN1(n951), .IN2(n849), .IN3(n935), .IN4(n941), .Q(n944) );
  INVX0 U879 ( .INP(n936), .ZN(n941) );
  NAND2X0 U880 ( .IN1(n799), .IN2(n797), .QN(n936) );
  NAND3X0 U881 ( .IN1(n952), .IN2(n953), .IN3(n849), .QN(n797) );
  AO21X1 U882 ( .IN1(n849), .IN2(n953), .IN3(n952), .Q(n799) );
  OA221X1 U883 ( .IN1(n954), .IN2(n955), .IN3(n956), .IN4(n794), .IN5(n957), 
        .Q(n914) );
  NAND4X0 U884 ( .IN1(n958), .IN2(n699), .IN3(n959), .IN4(n960), .QN(n957) );
  OA221X1 U885 ( .IN1(n714), .IN2(n705), .IN3(n713), .IN4(n712), .IN5(n961), 
        .Q(n960) );
  OA222X1 U886 ( .IN1(n704), .IN2(n708), .IN3(n711), .IN4(n767), .IN5(n707), 
        .IN6(n717), .Q(n961) );
  OA22X1 U887 ( .IN1(n716), .IN2(n757), .IN3(n702), .IN4(n732), .Q(n959) );
  NOR2X0 U888 ( .IN1(n694), .IN2(N33), .QN(n699) );
  XOR2X1 U889 ( .IN1(n962), .IN2(keyinput70), .Q(n958) );
  NAND2X0 U890 ( .IN1(n963), .IN2(N77), .QN(n962) );
  AOI221X1 U891 ( .IN1(n964), .IN2(n804), .IN3(n758), .IN4(n909), .IN5(n965), 
        .QN(n956) );
  AO221X1 U892 ( .IN1(N317), .IN2(n765), .IN3(N107), .IN4(n734), .IN5(n966), 
        .Q(n955) );
  AO21X1 U893 ( .IN1(N116), .IN2(n719), .IN3(n873), .Q(n966) );
  AO221X1 U894 ( .IN1(N303), .IN2(n833), .IN3(n963), .IN4(N97), .IN5(n967), 
        .Q(n954) );
  AO222X1 U895 ( .IN1(N294), .IN2(n816), .IN3(n968), .IN4(N311), .IN5(N283), 
        .IN6(n884), .Q(n967) );
  XOR2X1 U896 ( .IN1(n713), .IN2(keyinput63), .Q(n968) );
  OA21X1 U897 ( .IN1(n949), .IN2(n969), .IN3(n748), .Q(n913) );
  XOR2X1 U898 ( .IN1(keyinput40), .IN2(n798), .Q(n969) );
  XNOR2X1 U899 ( .IN1(n970), .IN2(n971), .Q(n949) );
  NOR2X0 U900 ( .IN1(n972), .IN2(n973), .QN(n971) );
  AO21X1 U901 ( .IN1(n974), .IN2(n975), .IN3(n976), .Q(N5002) );
  MUX21X1 U902 ( .IN1(n977), .IN2(n978), .S(n979), .Q(n976) );
  XOR2X1 U903 ( .IN1(n980), .IN2(keyinput43), .Q(n978) );
  NAND2X0 U904 ( .IN1(N116), .IN2(n981), .QN(n980) );
  NOR2X0 U905 ( .IN1(n974), .IN2(n982), .QN(n977) );
  XOR3X1 U906 ( .IN1(n983), .IN2(n856), .IN3(n777), .Q(n982) );
  AO221X1 U907 ( .IN1(n984), .IN2(n845), .IN3(n985), .IN4(n986), .IN5(n987), 
        .Q(n777) );
  XOR2X1 U908 ( .IN1(n988), .IN2(keyinput101), .Q(n987) );
  NAND4X0 U909 ( .IN1(n989), .IN2(n845), .IN3(n990), .IN4(n864), .QN(n988) );
  NOR2X0 U910 ( .IN1(n849), .IN2(n991), .QN(n984) );
  OA21X1 U911 ( .IN1(n738), .IN2(n866), .IN3(n850), .Q(n991) );
  AO21X1 U912 ( .IN1(n992), .IN2(n989), .IN3(n993), .Q(n856) );
  MUX21X1 U913 ( .IN1(n772), .IN2(n994), .S(n992), .Q(n983) );
  NAND2X0 U914 ( .IN1(n995), .IN2(n996), .QN(n994) );
  NAND3X0 U915 ( .IN1(n990), .IN2(n864), .IN3(n845), .QN(n996) );
  NAND2X0 U916 ( .IN1(n846), .IN2(n845), .QN(n772) );
  XOR2X1 U917 ( .IN1(n997), .IN2(n841), .Q(n845) );
  NAND2X0 U918 ( .IN1(keyinput97), .IN2(n840), .QN(n997) );
  AND2X1 U919 ( .IN1(n780), .IN2(n998), .Q(n840) );
  AND2X1 U920 ( .IN1(n865), .IN2(n864), .Q(n846) );
  INVX0 U921 ( .INP(n738), .ZN(n864) );
  XOR2X1 U922 ( .IN1(n999), .IN2(n1000), .Q(n738) );
  AND2X1 U923 ( .IN1(n1001), .IN2(n849), .Q(n1000) );
  AO22X1 U924 ( .IN1(N68), .IN2(n717), .IN3(n1002), .IN4(N77), .Q(n975) );
  MUX21X1 U925 ( .IN1(N68), .IN2(n1003), .S(N58), .Q(n1002) );
  NOR2X0 U926 ( .IN1(N68), .IN2(n717), .QN(n1003) );
  OAI22X1 U927 ( .IN1(n1004), .IN2(n1005), .IN3(n1006), .IN4(n1007), .QN(N4944) );
  AO21X1 U928 ( .IN1(n868), .IN2(n739), .IN3(n736), .Q(n1007) );
  INVX0 U929 ( .INP(n748), .ZN(n736) );
  AO222X1 U930 ( .IN1(n1008), .IN2(n1009), .IN3(n829), .IN4(n724), .IN5(n1010), 
        .IN6(n1011), .Q(n1006) );
  OA221X1 U931 ( .IN1(n707), .IN2(n728), .IN3(n711), .IN4(n727), .IN5(n1012), 
        .Q(n1011) );
  OA221X1 U932 ( .IN1(n758), .IN2(n1013), .IN3(n729), .IN4(n1014), .IN5(n1015), 
        .Q(n1012) );
  XOR2X1 U933 ( .IN1(keyinput62), .IN2(n719), .Q(n1014) );
  XOR2X1 U934 ( .IN1(keyinput61), .IN2(n963), .Q(n1013) );
  INVX0 U935 ( .INP(N283), .ZN(n727) );
  OA221X1 U936 ( .IN1(n713), .IN2(n730), .IN3(n704), .IN4(n725), .IN5(n1016), 
        .Q(n1010) );
  OA21X1 U937 ( .IN1(n714), .IN2(n811), .IN3(n813), .Q(n1016) );
  INVX0 U938 ( .INP(N311), .ZN(n811) );
  INVX0 U939 ( .INP(n696), .ZN(n829) );
  NAND2X0 U940 ( .IN1(n746), .IN2(n694), .QN(n696) );
  XOR2X1 U941 ( .IN1(n1017), .IN2(keyinput81), .Q(n1008) );
  NAND4X0 U942 ( .IN1(n1018), .IN2(n1019), .IN3(n1020), .IN4(n1021), .QN(n1017) );
  OA221X1 U943 ( .IN1(n704), .IN2(n712), .IN3(n707), .IN4(n767), .IN5(n1022), 
        .Q(n1021) );
  OA221X1 U944 ( .IN1(n1023), .IN2(n757), .IN3(n708), .IN4(n1024), .IN5(n1025), 
        .Q(n1022) );
  XOR2X1 U945 ( .IN1(keyinput57), .IN2(n816), .Q(n1024) );
  INVX0 U946 ( .INP(N150), .ZN(n708) );
  XOR2X1 U947 ( .IN1(n703), .IN2(keyinput56), .Q(n1023) );
  INVX0 U948 ( .INP(N143), .ZN(n712) );
  OA22X1 U949 ( .IN1(n713), .IN2(n705), .IN3(n714), .IN4(n709), .Q(n1020) );
  INVX0 U950 ( .INP(N132), .ZN(n709) );
  INVX0 U951 ( .INP(N137), .ZN(n705) );
  NAND2X0 U952 ( .IN1(N58), .IN2(n734), .QN(n1019) );
  XOR2X1 U953 ( .IN1(n1026), .IN2(keyinput69), .Q(n1018) );
  NAND2X0 U954 ( .IN1(n719), .IN2(N50), .QN(n1026) );
  INVX0 U955 ( .INP(n732), .ZN(n719) );
  OA22X1 U956 ( .IN1(n1027), .IN2(n1028), .IN3(n995), .IN4(n1029), .Q(n1005)
         );
  AOI21X1 U957 ( .IN1(n989), .IN2(n868), .IN3(n1028), .QN(n1029) );
  INVX0 U958 ( .INP(n867), .ZN(n989) );
  XNOR2X1 U959 ( .IN1(n1030), .IN2(keyinput105), .Q(n1028) );
  NAND2X0 U960 ( .IN1(n990), .IN2(n867), .QN(n1030) );
  INVX0 U961 ( .INP(n868), .ZN(n990) );
  AOI21X1 U962 ( .IN1(n867), .IN2(n995), .IN3(n865), .QN(n1027) );
  NOR2X0 U963 ( .IN1(n858), .IN2(n868), .QN(n865) );
  XOR2X1 U964 ( .IN1(n1031), .IN2(n1032), .Q(n868) );
  NAND2X0 U965 ( .IN1(n849), .IN2(n1033), .QN(n1031) );
  INVX0 U966 ( .INP(n858), .ZN(n995) );
  NOR2X0 U967 ( .IN1(n693), .IN2(n1034), .QN(n1004) );
  XOR2X1 U968 ( .IN1(keyinput50), .IN2(n689), .Q(n1034) );
  INVX0 U969 ( .INP(n686), .ZN(N4815) );
  MUX21X1 U970 ( .IN1(n1035), .IN2(n1036), .S(n748), .Q(n686) );
  NOR2X0 U971 ( .IN1(n693), .IN2(n689), .QN(n748) );
  NAND2X0 U972 ( .IN1(N1), .IN2(n1037), .QN(n693) );
  NAND3X0 U973 ( .IN1(N13), .IN2(n1038), .IN3(N45), .QN(n1037) );
  AO221X1 U974 ( .IN1(n1039), .IN2(n1009), .IN3(n1040), .IN4(n798), .IN5(n1041), .Q(n1036) );
  AO22X1 U975 ( .IN1(n1042), .IN2(n1043), .IN3(n1044), .IN4(n1045), .Q(n1041)
         );
  AO222X1 U976 ( .IN1(n909), .IN2(n728), .IN3(n1046), .IN4(n804), .IN5(n965), 
        .IN6(N1947), .Q(n1045) );
  INVX0 U977 ( .INP(n803), .ZN(n965) );
  INVX0 U978 ( .INP(n901), .ZN(n804) );
  MUX21X1 U979 ( .IN1(n1047), .IN2(n1048), .S(n904), .Q(n1046) );
  XOR2X1 U980 ( .IN1(N45), .IN2(keyinput6), .Q(n904) );
  INVX0 U981 ( .INP(n800), .ZN(n909) );
  NAND2X0 U982 ( .IN1(n803), .IN2(n901), .QN(n800) );
  NAND2X0 U983 ( .IN1(N33), .IN2(n1049), .QN(n901) );
  NAND2X0 U984 ( .IN1(n1049), .IN2(n1025), .QN(n803) );
  XOR2X1 U985 ( .IN1(n1050), .IN2(keyinput10), .Q(n1049) );
  INVX0 U986 ( .INP(n794), .ZN(n1044) );
  NAND2X0 U987 ( .IN1(n876), .IN2(n694), .QN(n794) );
  INVX0 U988 ( .INP(n1009), .ZN(n694) );
  OA221X1 U989 ( .IN1(n732), .IN2(n730), .IN3(n716), .IN4(n725), .IN5(n1051), 
        .Q(n1043) );
  AOI222X1 U990 ( .IN1(N329), .IN2(n765), .IN3(N311), .IN4(n884), .IN5(N283), 
        .IN6(n963), .QN(n1051) );
  INVX0 U991 ( .INP(n703), .ZN(n963) );
  INVX0 U992 ( .INP(n707), .ZN(n884) );
  INVX0 U993 ( .INP(n714), .ZN(n765) );
  INVX0 U994 ( .INP(N294), .ZN(n725) );
  INVX0 U995 ( .INP(N303), .ZN(n730) );
  OA221X1 U996 ( .IN1(n704), .IN2(n809), .IN3(n711), .IN4(n812), .IN5(n1052), 
        .Q(n1042) );
  OA21X1 U997 ( .IN1(n713), .IN2(n892), .IN3(n813), .Q(n1052) );
  INVX0 U998 ( .INP(n873), .ZN(n813) );
  NAND2X0 U999 ( .IN1(N33), .IN2(n1009), .QN(n873) );
  INVX0 U1000 ( .INP(N326), .ZN(n892) );
  INVX0 U1001 ( .INP(N317), .ZN(n812) );
  INVX0 U1002 ( .INP(N322), .ZN(n809) );
  INVX0 U1003 ( .INP(n876), .ZN(n798) );
  NAND2X0 U1004 ( .IN1(n739), .IN2(n1038), .QN(n876) );
  INVX0 U1005 ( .INP(n746), .ZN(n739) );
  NAND2X0 U1006 ( .IN1(n1053), .IN2(n1025), .QN(n746) );
  XOR2X1 U1007 ( .IN1(keyinput3), .IN2(n1054), .Q(n1053) );
  XOR2X1 U1008 ( .IN1(n1055), .IN2(n1056), .Q(n1040) );
  OA21X1 U1009 ( .IN1(n1038), .IN2(N169), .IN3(n1057), .Q(n1009) );
  XOR2X1 U1010 ( .IN1(n1058), .IN2(keyinput82), .Q(n1039) );
  NAND4X0 U1011 ( .IN1(n1059), .IN2(n1060), .IN3(n1061), .IN4(n1062), .QN(
        n1058) );
  OA221X1 U1012 ( .IN1(n732), .IN2(n758), .IN3(n714), .IN4(n767), .IN5(n1063), 
        .Q(n1062) );
  OA22X1 U1013 ( .IN1(n713), .IN2(n717), .IN3(n703), .IN4(n729), .Q(n1063) );
  NAND2X0 U1014 ( .IN1(n1064), .IN2(n1065), .QN(n703) );
  XOR2X1 U1015 ( .IN1(n1066), .IN2(keyinput39), .Q(n713) );
  NAND2X0 U1016 ( .IN1(n1067), .IN2(N200), .QN(n1066) );
  NAND2X0 U1017 ( .IN1(n1065), .IN2(n1068), .QN(n714) );
  NAND2X0 U1018 ( .IN1(n1064), .IN2(n1069), .QN(n732) );
  AND3X1 U1019 ( .IN1(N20), .IN2(n1070), .IN3(N200), .Q(n1064) );
  OA22X1 U1020 ( .IN1(n707), .IN2(n724), .IN3(n704), .IN4(n702), .Q(n1061) );
  INVX0 U1021 ( .INP(n833), .ZN(n704) );
  XOR2X1 U1022 ( .IN1(n1071), .IN2(keyinput38), .Q(n833) );
  NAND2X0 U1023 ( .IN1(n1067), .IN2(n1072), .QN(n1071) );
  NOR2X0 U1024 ( .IN1(n1073), .IN2(n1065), .QN(n1067) );
  NAND3X0 U1025 ( .IN1(n1074), .IN2(n1072), .IN3(n1065), .QN(n707) );
  NAND2X0 U1026 ( .IN1(N68), .IN2(n816), .QN(n1060) );
  INVX0 U1027 ( .INP(n711), .ZN(n816) );
  NAND3X0 U1028 ( .IN1(n1074), .IN2(N200), .IN3(n1065), .QN(n711) );
  INVX0 U1029 ( .INP(n1069), .ZN(n1065) );
  AND2X1 U1030 ( .IN1(n1025), .IN2(n1015), .Q(n1059) );
  NAND2X0 U1031 ( .IN1(N97), .IN2(n734), .QN(n1015) );
  INVX0 U1032 ( .INP(n716), .ZN(n734) );
  NAND2X0 U1033 ( .IN1(n1068), .IN2(n1069), .QN(n716) );
  NAND2X0 U1034 ( .IN1(n1075), .IN2(n1076), .QN(n1069) );
  XOR2X1 U1035 ( .IN1(keyinput7), .IN2(N20), .Q(n1075) );
  OA21X1 U1036 ( .IN1(n1072), .IN2(n1038), .IN3(n1070), .Q(n1068) );
  XNOR2X1 U1037 ( .IN1(n1073), .IN2(keyinput13), .Q(n1070) );
  INVX0 U1038 ( .INP(n1074), .ZN(n1073) );
  NOR2X0 U1039 ( .IN1(n1077), .IN2(n1038), .QN(n1074) );
  AO21X1 U1040 ( .IN1(n1078), .IN2(n1079), .IN3(n1080), .Q(n1035) );
  AO21X1 U1041 ( .IN1(n923), .IN2(n1081), .IN3(n1082), .Q(N4667) );
  MUX21X1 U1042 ( .IN1(n1083), .IN2(n1084), .S(n689), .Q(n1082) );
  INVX0 U1043 ( .INP(n869), .ZN(n689) );
  NAND2X0 U1044 ( .IN1(n1050), .IN2(n1085), .QN(n869) );
  INVX0 U1045 ( .INP(n1048), .ZN(n1084) );
  NOR2X0 U1046 ( .IN1(n1081), .IN2(n908), .QN(n1083) );
  NAND4X0 U1047 ( .IN1(n729), .IN2(n728), .IN3(n758), .IN4(n731), .QN(n908) );
  NAND2X0 U1048 ( .IN1(n858), .IN2(n867), .QN(n923) );
  NAND2X0 U1049 ( .IN1(n1086), .IN2(n973), .QN(n867) );
  AO21X1 U1050 ( .IN1(n1087), .IN2(n1088), .IN3(n1079), .Q(n858) );
  INVX0 U1051 ( .INP(N330), .ZN(n1079) );
  NAND2X0 U1052 ( .IN1(n1089), .IN2(n973), .QN(n1088) );
  XNOR2X1 U1053 ( .IN1(keyinput83), .IN2(n1090), .Q(n1087) );
  NOR2X0 U1054 ( .IN1(n973), .IN2(n1091), .QN(n1090) );
  MUX21X1 U1055 ( .IN1(n1092), .IN2(n1093), .S(n1094), .Q(n1091) );
  NAND3X0 U1056 ( .IN1(n1095), .IN2(n1096), .IN3(n1097), .QN(n1093) );
  INVX0 U1057 ( .INP(n1098), .ZN(n1096) );
  NAND4X0 U1058 ( .IN1(n1099), .IN2(n1098), .IN3(n1100), .IN4(n1101), .QN(
        n1092) );
  XNOR2X1 U1059 ( .IN1(N179), .IN2(keyinput15), .Q(n1099) );
  NAND2X0 U1060 ( .IN1(n935), .IN2(n930), .QN(N4589) );
  NAND2X0 U1061 ( .IN1(n1080), .IN2(n875), .QN(n930) );
  INVX0 U1062 ( .INP(n910), .ZN(n1080) );
  NAND2X0 U1063 ( .IN1(N330), .IN2(n943), .QN(n910) );
  INVX0 U1064 ( .INP(n1078), .ZN(n943) );
  XOR2X1 U1065 ( .IN1(n1102), .IN2(n1103), .Q(n1078) );
  NOR2X0 U1066 ( .IN1(keyinput95), .IN2(n1055), .QN(n1103) );
  NAND2X0 U1067 ( .IN1(n849), .IN2(n1104), .QN(n1055) );
  AOI21X1 U1068 ( .IN1(n929), .IN2(n875), .IN3(n1105), .QN(n935) );
  XOR2X1 U1069 ( .IN1(n1106), .IN2(keyinput93), .Q(n1105) );
  OR2X1 U1070 ( .IN1(n1107), .IN2(n849), .Q(n1106) );
  XOR3X1 U1071 ( .IN1(keyinput67), .IN2(n1108), .IN3(n1109), .Q(n875) );
  AND2X1 U1072 ( .IN1(n1110), .IN2(n849), .Q(n1108) );
  NOR2X0 U1073 ( .IN1(n1111), .IN2(n849), .QN(n929) );
  INVX0 U1074 ( .INP(n973), .ZN(n849) );
  NAND2X0 U1075 ( .IN1(N343), .IN2(n780), .QN(n973) );
  INVX0 U1076 ( .INP(n986), .ZN(n780) );
  NAND3X0 U1077 ( .IN1(N213), .IN2(n1038), .IN3(n1112), .QN(n986) );
  MUX21X1 U1078 ( .IN1(n1113), .IN2(n1057), .S(keyinput1), .Q(n1112) );
  NOR2X0 U1079 ( .IN1(N1), .IN2(n1054), .QN(n1113) );
  AO21X1 U1080 ( .IN1(n992), .IN2(n1086), .IN3(n993), .Q(N4145) );
  OAI21X1 U1081 ( .IN1(n1114), .IN2(n779), .IN3(n1115), .QN(n993) );
  OA21X1 U1082 ( .IN1(n1116), .IN2(n841), .IN3(n1117), .Q(n1114) );
  OA21X1 U1083 ( .IN1(n999), .IN2(n866), .IN3(n850), .Q(n1116) );
  XNOR2X1 U1084 ( .IN1(n1118), .IN2(keyinput87), .Q(n866) );
  INVX0 U1085 ( .INP(n1119), .ZN(n999) );
  XOR2X1 U1086 ( .IN1(keyinput94), .IN2(n1120), .Q(n1086) );
  OA21X1 U1087 ( .IN1(n1121), .IN2(n970), .IN3(n1122), .Q(n1120) );
  XNOR2X1 U1088 ( .IN1(keyinput91), .IN2(n1123), .Q(n1122) );
  OA21X1 U1089 ( .IN1(n1124), .IN2(n952), .IN3(n951), .Q(n1121) );
  OA21X1 U1090 ( .IN1(n1109), .IN2(n1111), .IN3(n1107), .Q(n1124) );
  AND2X1 U1091 ( .IN1(n1089), .IN2(n992), .Q(N4028) );
  INVX0 U1092 ( .INP(n859), .ZN(n992) );
  NAND4X0 U1093 ( .IN1(n1125), .IN2(n1032), .IN3(n1119), .IN4(n1126), .QN(n859) );
  INVX0 U1094 ( .INP(n779), .ZN(n1126) );
  XNOR2X1 U1095 ( .IN1(keyinput89), .IN2(n1127), .Q(n779) );
  OA21X1 U1096 ( .IN1(n781), .IN2(n1128), .IN3(n1115), .Q(n1127) );
  AND2X1 U1097 ( .IN1(n1129), .IN2(n1130), .Q(n1115) );
  NAND3X0 U1098 ( .IN1(n1131), .IN2(n781), .IN3(N169), .QN(n1130) );
  XNOR2X1 U1099 ( .IN1(n1132), .IN2(keyinput77), .Q(n1129) );
  NAND3X0 U1100 ( .IN1(N179), .IN2(n781), .IN3(n1133), .QN(n1132) );
  MUX21X1 U1101 ( .IN1(N200), .IN2(N190), .S(n1133), .Q(n1128) );
  INVX0 U1102 ( .INP(n1131), .ZN(n1133) );
  AO221X1 U1103 ( .IN1(n1134), .IN2(n1135), .IN3(n1136), .IN4(N226), .IN5(
        n1137), .Q(n1131) );
  AO222X1 U1104 ( .IN1(N222), .IN2(n1138), .IN3(N223), .IN4(n1139), .IN5(N33), 
        .IN6(N77), .Q(n1135) );
  AO21X1 U1105 ( .IN1(n1140), .IN2(n1141), .IN3(n1142), .Q(n781) );
  MUX21X1 U1106 ( .IN1(n1143), .IN2(n1144), .S(N50), .Q(n1142) );
  AO221X1 U1107 ( .IN1(n1145), .IN2(n1146), .IN3(N150), .IN4(n1147), .IN5(
        n1148), .Q(n1140) );
  XOR2X1 U1108 ( .IN1(keyinput21), .IN2(n1149), .Q(n1148) );
  NOR2X0 U1109 ( .IN1(n702), .IN2(n1150), .QN(n1149) );
  XOR2X1 U1110 ( .IN1(n1038), .IN2(keyinput11), .Q(n1145) );
  OA21X1 U1111 ( .IN1(n1151), .IN2(n1001), .IN3(n850), .Q(n1119) );
  NAND2X0 U1112 ( .IN1(n1152), .IN2(n1001), .QN(n850) );
  MUX21X1 U1113 ( .IN1(N169), .IN2(N179), .S(n1153), .Q(n1152) );
  AO21X1 U1114 ( .IN1(n1154), .IN2(n1141), .IN3(n1155), .Q(n1001) );
  MUX21X1 U1115 ( .IN1(n1143), .IN2(n1144), .S(N68), .Q(n1155) );
  AO222X1 U1116 ( .IN1(n1156), .IN2(N77), .IN3(N50), .IN4(n1157), .IN5(N20), 
        .IN6(n757), .Q(n1154) );
  XOR2X1 U1117 ( .IN1(keyinput18), .IN2(n1147), .Q(n1157) );
  MUX21X1 U1118 ( .IN1(N200), .IN2(N190), .S(n1153), .Q(n1151) );
  AOI221X1 U1119 ( .IN1(n1134), .IN2(n1158), .IN3(n1136), .IN4(N238), .IN5(
        n1137), .QN(n1153) );
  AO222X1 U1120 ( .IN1(N232), .IN2(n1139), .IN3(N97), .IN4(n1159), .IN5(N226), 
        .IN6(n1138), .Q(n1158) );
  XOR2X1 U1121 ( .IN1(keyinput23), .IN2(N33), .Q(n1159) );
  OA21X1 U1122 ( .IN1(n1160), .IN2(n1033), .IN3(n1118), .Q(n1032) );
  NAND3X0 U1123 ( .IN1(n1161), .IN2(n1033), .IN3(n1162), .QN(n1118) );
  MUX21X1 U1124 ( .IN1(n1163), .IN2(n1164), .S(keyinput65), .Q(n1162) );
  NAND2X0 U1125 ( .IN1(n1163), .IN2(n1165), .QN(n1164) );
  INVX0 U1126 ( .INP(N169), .ZN(n1165) );
  AO21X1 U1127 ( .IN1(N169), .IN2(n1163), .IN3(N179), .Q(n1161) );
  AO21X1 U1128 ( .IN1(n1166), .IN2(n1141), .IN3(n1167), .Q(n1033) );
  MUX21X1 U1129 ( .IN1(n1143), .IN2(n1168), .S(N77), .Q(n1167) );
  MUX21X1 U1130 ( .IN1(n1144), .IN2(n1169), .S(keyinput25), .Q(n1168) );
  NOR2X0 U1131 ( .IN1(n1170), .IN2(n1171), .QN(n1169) );
  XOR2X1 U1132 ( .IN1(keyinput28), .IN2(n1172), .Q(n1166) );
  OA221X1 U1133 ( .IN1(n702), .IN2(n1173), .IN3(n1038), .IN4(n724), .IN5(n1174), .Q(n1172) );
  XOR2X1 U1134 ( .IN1(keyinput22), .IN2(n1175), .Q(n1174) );
  NOR2X0 U1135 ( .IN1(n758), .IN2(n1150), .QN(n1175) );
  INVX0 U1136 ( .INP(N77), .ZN(n724) );
  OA22X1 U1137 ( .IN1(n1176), .IN2(n1163), .IN3(N200), .IN4(n1177), .Q(n1160)
         );
  AOI21X1 U1138 ( .IN1(n1163), .IN2(keyinput65), .IN3(n1076), .QN(n1177) );
  AO221X1 U1139 ( .IN1(n1134), .IN2(n1178), .IN3(n1136), .IN4(N244), .IN5(
        n1137), .Q(n1163) );
  AO222X1 U1140 ( .IN1(N232), .IN2(n1138), .IN3(N238), .IN4(n1139), .IN5(N33), 
        .IN6(N107), .Q(n1178) );
  AND2X1 U1141 ( .IN1(N190), .IN2(keyinput65), .Q(n1176) );
  INVX0 U1142 ( .INP(n841), .ZN(n1125) );
  NAND2X0 U1143 ( .IN1(n1179), .IN2(n1117), .QN(n841) );
  INVX0 U1144 ( .INP(n985), .ZN(n1117) );
  NAND2X0 U1145 ( .IN1(n1180), .IN2(n1181), .QN(n985) );
  NAND3X0 U1146 ( .IN1(n998), .IN2(n1182), .IN3(N169), .QN(n1181) );
  XOR2X1 U1147 ( .IN1(n1183), .IN2(keyinput86), .Q(n1180) );
  NAND3X0 U1148 ( .IN1(N179), .IN2(n998), .IN3(n1184), .QN(n1183) );
  XOR2X1 U1149 ( .IN1(n1185), .IN2(keyinput78), .Q(n998) );
  XOR2X1 U1150 ( .IN1(n1186), .IN2(keyinput90), .Q(n1179) );
  NAND2X0 U1151 ( .IN1(n1187), .IN2(n1185), .QN(n1186) );
  AOI21X1 U1152 ( .IN1(n1141), .IN2(n1188), .IN3(n1189), .QN(n1185) );
  MUX21X1 U1153 ( .IN1(n1143), .IN2(n1144), .S(N58), .Q(n1189) );
  NOR2X0 U1154 ( .IN1(n1190), .IN2(n1171), .QN(n1144) );
  NOR2X0 U1155 ( .IN1(n1038), .IN2(N1), .QN(n1171) );
  INVX0 U1156 ( .INP(n1170), .ZN(n1190) );
  OAI21X1 U1157 ( .IN1(n767), .IN2(n1173), .IN3(n1191), .QN(n1188) );
  MUX21X1 U1158 ( .IN1(n1192), .IN2(n1193), .S(N68), .Q(n1191) );
  OA21X1 U1159 ( .IN1(n1038), .IN2(n702), .IN3(n1150), .Q(n1193) );
  NAND2X0 U1160 ( .IN1(N20), .IN2(n702), .QN(n1192) );
  INVX0 U1161 ( .INP(N159), .ZN(n767) );
  MUX21X1 U1162 ( .IN1(n1072), .IN2(n1076), .S(n1184), .Q(n1187) );
  INVX0 U1163 ( .INP(n1182), .ZN(n1184) );
  AO221X1 U1164 ( .IN1(n1194), .IN2(n1134), .IN3(n1136), .IN4(N232), .IN5(
        n1137), .Q(n1182) );
  AND3X1 U1165 ( .IN1(N274), .IN2(n1195), .IN3(n1196), .Q(n1137) );
  NOR2X0 U1166 ( .IN1(n1196), .IN2(n1134), .QN(n1136) );
  XOR2X1 U1167 ( .IN1(n1197), .IN2(keyinput9), .Q(n1196) );
  NAND2X0 U1168 ( .IN1(n1198), .IN2(n1199), .QN(n1197) );
  XOR2X1 U1169 ( .IN1(keyinput5), .IN2(n1200), .Q(n1198) );
  NOR2X0 U1170 ( .IN1(N41), .IN2(N45), .QN(n1200) );
  XOR2X1 U1171 ( .IN1(n1201), .IN2(keyinput41), .Q(n1194) );
  AO221X1 U1172 ( .IN1(n1202), .IN2(N223), .IN3(N33), .IN4(N87), .IN5(n1203), 
        .Q(n1201) );
  XOR2X1 U1173 ( .IN1(n1204), .IN2(keyinput29), .Q(n1203) );
  NAND2X0 U1174 ( .IN1(N226), .IN2(n1139), .QN(n1204) );
  XNOR2X1 U1175 ( .IN1(n1138), .IN2(keyinput14), .Q(n1202) );
  NOR4X0 U1176 ( .IN1(n970), .IN2(n952), .IN3(n1109), .IN4(n1102), .QN(n1089)
         );
  INVX0 U1177 ( .INP(n1056), .ZN(n1102) );
  OA21X1 U1178 ( .IN1(n1205), .IN2(n1104), .IN3(n1111), .Q(n1056) );
  NAND2X0 U1179 ( .IN1(n1206), .IN2(n1104), .QN(n1111) );
  MUX21X1 U1180 ( .IN1(N169), .IN2(N179), .S(n1094), .Q(n1206) );
  AO21X1 U1181 ( .IN1(n1207), .IN2(n1141), .IN3(n1208), .Q(n1104) );
  MUX21X1 U1182 ( .IN1(n1143), .IN2(n1209), .S(N116), .Q(n1208) );
  AO22X1 U1183 ( .IN1(N283), .IN2(n1156), .IN3(n1147), .IN4(N97), .Q(n1207) );
  MUX21X1 U1184 ( .IN1(N200), .IN2(N190), .S(n1094), .Q(n1205) );
  AOI221X1 U1185 ( .IN1(N270), .IN2(n1210), .IN3(n1134), .IN4(n1211), .IN5(
        n1212), .QN(n1094) );
  AO221X1 U1186 ( .IN1(N264), .IN2(n1139), .IN3(N303), .IN4(N33), .IN5(n1213), 
        .Q(n1211) );
  XOR2X1 U1187 ( .IN1(n1214), .IN2(keyinput19), .Q(n1213) );
  NAND2X0 U1188 ( .IN1(N257), .IN2(n1138), .QN(n1214) );
  NAND2X0 U1189 ( .IN1(n1215), .IN2(n1216), .QN(n1109) );
  AO221X1 U1190 ( .IN1(n1217), .IN2(N190), .IN3(n1098), .IN4(N200), .IN5(n1110), .Q(n1216) );
  XOR2X1 U1191 ( .IN1(n1107), .IN2(keyinput88), .Q(n1215) );
  NAND2X0 U1192 ( .IN1(n1218), .IN2(n1110), .QN(n1107) );
  AO21X1 U1193 ( .IN1(n1219), .IN2(n1141), .IN3(n1220), .Q(n1110) );
  MUX21X1 U1194 ( .IN1(n1143), .IN2(n1221), .S(N107), .Q(n1220) );
  AO222X1 U1195 ( .IN1(n1147), .IN2(N87), .IN3(n1222), .IN4(n729), .IN5(N116), 
        .IN6(n1156), .Q(n1219) );
  XOR2X1 U1196 ( .IN1(n1038), .IN2(keyinput12), .Q(n1222) );
  AO22X1 U1197 ( .IN1(N169), .IN2(n1098), .IN3(n1217), .IN4(N179), .Q(n1218)
         );
  XOR2X1 U1198 ( .IN1(n1098), .IN2(keyinput66), .Q(n1217) );
  XOR2X1 U1199 ( .IN1(n1223), .IN2(keyinput48), .Q(n1098) );
  AO221X1 U1200 ( .IN1(N264), .IN2(n1210), .IN3(n1134), .IN4(n1224), .IN5(
        n1212), .Q(n1223) );
  INVX0 U1201 ( .INP(n1225), .ZN(n1212) );
  AO222X1 U1202 ( .IN1(N250), .IN2(n1138), .IN3(N257), .IN4(n1226), .IN5(N294), 
        .IN6(N33), .Q(n1224) );
  XOR2X1 U1203 ( .IN1(keyinput24), .IN2(n1139), .Q(n1226) );
  OAI21X1 U1204 ( .IN1(n1227), .IN2(n953), .IN3(n951), .QN(n952) );
  NAND2X0 U1205 ( .IN1(n1228), .IN2(n953), .QN(n951) );
  MUX21X1 U1206 ( .IN1(N169), .IN2(N179), .S(n1097), .Q(n1228) );
  INVX0 U1207 ( .INP(n1100), .ZN(n1097) );
  AO221X1 U1208 ( .IN1(n1229), .IN2(n1141), .IN3(n1143), .IN4(n731), .IN5(
        n1230), .Q(n953) );
  XOR2X1 U1209 ( .IN1(keyinput31), .IN2(n1231), .Q(n1230) );
  AND2X1 U1210 ( .IN1(N97), .IN2(n1221), .Q(n1231) );
  AO222X1 U1211 ( .IN1(n1147), .IN2(N77), .IN3(N20), .IN4(n1232), .IN5(n1156), 
        .IN6(N107), .Q(n1229) );
  INVX0 U1212 ( .INP(n1150), .ZN(n1156) );
  XOR2X1 U1213 ( .IN1(keyinput36), .IN2(n981), .Q(n1232) );
  XOR2X1 U1214 ( .IN1(N97), .IN2(N107), .Q(n981) );
  MUX21X1 U1215 ( .IN1(N190), .IN2(N200), .S(n1100), .Q(n1227) );
  NAND3X0 U1216 ( .IN1(n1233), .IN2(n1225), .IN3(n1234), .QN(n1100) );
  XOR2X1 U1217 ( .IN1(keyinput45), .IN2(n1235), .Q(n1234) );
  NOR2X0 U1218 ( .IN1(n1236), .IN2(n1195), .QN(n1235) );
  INVX0 U1219 ( .INP(n1134), .ZN(n1195) );
  XOR2X1 U1220 ( .IN1(n1237), .IN2(keyinput42), .Q(n1236) );
  AO222X1 U1221 ( .IN1(N244), .IN2(n1138), .IN3(N250), .IN4(n1139), .IN5(N283), 
        .IN6(N33), .Q(n1237) );
  NAND3X0 U1222 ( .IN1(n1238), .IN2(n1239), .IN3(N274), .QN(n1225) );
  INVX0 U1223 ( .INP(n1240), .ZN(n1238) );
  NAND2X0 U1224 ( .IN1(N257), .IN2(n1210), .QN(n1233) );
  AND2X1 U1225 ( .IN1(n1239), .IN2(n1240), .Q(n1210) );
  NAND3X0 U1226 ( .IN1(n1199), .IN2(n1085), .IN3(N45), .QN(n1240) );
  XOR2X1 U1227 ( .IN1(N1), .IN2(keyinput2), .Q(n1199) );
  AO21X1 U1228 ( .IN1(n1241), .IN2(n972), .IN3(n1123), .Q(n970) );
  NAND2X0 U1229 ( .IN1(n1242), .IN2(n1243), .QN(n1123) );
  NAND3X0 U1230 ( .IN1(n1244), .IN2(n1101), .IN3(N169), .QN(n1243) );
  XOR2X1 U1231 ( .IN1(n1245), .IN2(keyinput79), .Q(n1242) );
  NAND2X0 U1232 ( .IN1(n1095), .IN2(n1244), .QN(n1245) );
  NOR2X0 U1233 ( .IN1(n1101), .IN2(n1077), .QN(n1095) );
  INVX0 U1234 ( .INP(N179), .ZN(n1077) );
  INVX0 U1235 ( .INP(n1244), .ZN(n972) );
  AO221X1 U1236 ( .IN1(n1246), .IN2(n1141), .IN3(N87), .IN4(n1209), .IN5(n1247), .Q(n1244) );
  XOR2X1 U1237 ( .IN1(keyinput26), .IN2(n1248), .Q(n1247) );
  NOR2X0 U1238 ( .IN1(N87), .IN2(n1249), .QN(n1248) );
  AO21X1 U1239 ( .IN1(N20), .IN2(n1141), .IN3(n1221), .Q(n1209) );
  OA21X1 U1240 ( .IN1(n1025), .IN2(N1), .IN3(n1170), .Q(n1221) );
  NOR2X0 U1241 ( .IN1(n1141), .IN2(n1143), .QN(n1170) );
  INVX0 U1242 ( .INP(n1249), .ZN(n1143) );
  NAND2X0 U1243 ( .IN1(n1250), .IN2(n1081), .QN(n1249) );
  XOR3X1 U1244 ( .IN1(keyinput8), .IN2(keyinput4), .IN3(n1251), .Q(n1250) );
  NOR2X0 U1245 ( .IN1(n1054), .IN2(n1038), .QN(n1251) );
  INVX0 U1246 ( .INP(N13), .ZN(n1054) );
  NAND2X0 U1247 ( .IN1(n1252), .IN2(n1253), .QN(n1141) );
  NAND3X0 U1248 ( .IN1(N20), .IN2(N1), .IN3(N33), .QN(n1253) );
  AO21X1 U1249 ( .IN1(N107), .IN2(N20), .IN3(n1254), .Q(n1246) );
  MUX21X1 U1250 ( .IN1(N97), .IN2(N68), .S(n1147), .Q(n1254) );
  INVX0 U1251 ( .INP(n1173), .ZN(n1147) );
  NAND2X0 U1252 ( .IN1(n1038), .IN2(n1150), .QN(n1173) );
  NAND2X0 U1253 ( .IN1(N33), .IN2(n1038), .QN(n1150) );
  INVX0 U1254 ( .INP(N20), .ZN(n1038) );
  MUX21X1 U1255 ( .IN1(n1076), .IN2(n1072), .S(n1101), .Q(n1241) );
  AO22X1 U1256 ( .IN1(n1134), .IN2(n1255), .IN3(n1256), .IN4(n1239), .Q(n1101)
         );
  XOR2X1 U1257 ( .IN1(n1134), .IN2(keyinput30), .Q(n1239) );
  MUX21X1 U1258 ( .IN1(N250), .IN2(N274), .S(n1257), .Q(n1256) );
  NOR2X0 U1259 ( .IN1(n1258), .IN2(n1259), .QN(n1257) );
  XOR2X1 U1260 ( .IN1(keyinput1), .IN2(N1), .Q(n1259) );
  INVX0 U1261 ( .INP(N45), .ZN(n1258) );
  AO222X1 U1262 ( .IN1(N238), .IN2(n1138), .IN3(N244), .IN4(n1139), .IN5(N116), 
        .IN6(N33), .Q(n1255) );
  NOR2X0 U1263 ( .IN1(n1138), .IN2(N33), .QN(n1139) );
  NOR2X0 U1264 ( .IN1(N349), .IN2(N33), .QN(n1138) );
  OA21X1 U1265 ( .IN1(n1085), .IN2(n1025), .IN3(n1057), .Q(n1134) );
  INVX0 U1266 ( .INP(N33), .ZN(n1025) );
  INVX0 U1267 ( .INP(N41), .ZN(n1085) );
  INVX0 U1268 ( .INP(N200), .ZN(n1072) );
  INVX0 U1269 ( .INP(N190), .ZN(n1076) );
  XOR2X1 U1270 ( .IN1(n1047), .IN2(n801), .Q(N3987) );
  XOR3X1 U1271 ( .IN1(n729), .IN2(n1260), .IN3(n1261), .Q(n801) );
  XOR2X1 U1272 ( .IN1(n728), .IN2(N87), .Q(n1261) );
  INVX0 U1273 ( .INP(N116), .ZN(n728) );
  NOR2X0 U1274 ( .IN1(N97), .IN2(keyinput27), .QN(n1260) );
  XOR3X1 U1275 ( .IN1(N50), .IN2(n1262), .IN3(n1263), .Q(n1047) );
  NAND2X0 U1276 ( .IN1(keyinput17), .IN2(n830), .QN(n1263) );
  XOR2X1 U1277 ( .IN1(N77), .IN2(N68), .Q(n1262) );
  AO22X1 U1278 ( .IN1(n1264), .IN2(n1265), .IN3(keyinput92), .IN4(n1266), .Q(
        N3833) );
  NAND2X0 U1279 ( .IN1(keyinput84), .IN2(n1265), .QN(n1266) );
  OR2X1 U1280 ( .IN1(n1267), .IN2(n964), .Q(n1265) );
  NAND3X0 U1281 ( .IN1(n1268), .IN2(n1267), .IN3(n964), .QN(n1264) );
  XNOR3X1 U1282 ( .IN1(N257), .IN2(N250), .IN3(n1269), .Q(n964) );
  XNOR2X1 U1283 ( .IN1(N270), .IN2(N264), .Q(n1269) );
  AO21X1 U1284 ( .IN1(keyinput46), .IN2(n1270), .IN3(n1271), .Q(n1267) );
  MUX21X1 U1285 ( .IN1(n1272), .IN2(n1273), .S(n907), .Q(n1271) );
  XOR2X1 U1286 ( .IN1(N238), .IN2(N244), .Q(n907) );
  NOR2X0 U1287 ( .IN1(keyinput46), .IN2(n1272), .QN(n1273) );
  NAND2X0 U1288 ( .IN1(keyinput47), .IN2(n906), .QN(n1272) );
  INVX0 U1289 ( .INP(n1270), .ZN(n906) );
  XOR3X1 U1290 ( .IN1(keyinput20), .IN2(N232), .IN3(N226), .Q(n1270) );
  NAND2X0 U1291 ( .IN1(keyinput84), .IN2(n1274), .QN(n1268) );
  INVX0 U1292 ( .INP(keyinput92), .ZN(n1274) );
  NOR2X0 U1293 ( .IN1(N77), .IN2(n1146), .QN(N1713) );
  NAND3X0 U1294 ( .IN1(n702), .IN2(n757), .IN3(n717), .QN(n1146) );
  INVX0 U1295 ( .INP(N58), .ZN(n702) );
  AOI221X1 U1296 ( .IN1(n1275), .IN2(N250), .IN3(n1276), .IN4(n1277), .IN5(
        n1278), .QN(N3195) );
  XOR2X1 U1297 ( .IN1(keyinput44), .IN2(n1279), .Q(n1278) );
  NOR2X0 U1298 ( .IN1(n1048), .IN2(n1280), .QN(n1279) );
  AO21X1 U1299 ( .IN1(n830), .IN2(n757), .IN3(n717), .Q(n1048) );
  INVX0 U1300 ( .INP(N50), .ZN(n717) );
  INVX0 U1301 ( .INP(N68), .ZN(n757) );
  XOR2X1 U1302 ( .IN1(N58), .IN2(keyinput0), .Q(n830) );
  NAND4X0 U1303 ( .IN1(n1281), .IN2(n1282), .IN3(n1283), .IN4(n1284), .QN(
        n1277) );
  AOI22X1 U1304 ( .IN1(N107), .IN2(N264), .IN3(N116), .IN4(N270), .QN(n1284)
         );
  AOI22X1 U1305 ( .IN1(N50), .IN2(N226), .IN3(N58), .IN4(N232), .QN(n1283) );
  AOI22X1 U1306 ( .IN1(N68), .IN2(N238), .IN3(N77), .IN4(N244), .QN(n1282) );
  AOI22X1 U1307 ( .IN1(N87), .IN2(N250), .IN3(N97), .IN4(N257), .QN(n1281) );
  XOR2X1 U1308 ( .IN1(keyinput37), .IN2(n1285), .Q(n1276) );
  NOR2X0 U1309 ( .IN1(n979), .IN2(n1050), .QN(n1285) );
  INVX0 U1310 ( .INP(n1280), .ZN(n979) );
  NAND2X0 U1311 ( .IN1(N20), .IN2(n1057), .QN(n1280) );
  OA21X1 U1312 ( .IN1(N264), .IN2(N257), .IN3(n1050), .Q(n1275) );
  AND2X1 U1313 ( .IN1(N20), .IN2(n974), .Q(n1050) );
  MUX21X1 U1314 ( .IN1(n1286), .IN2(n1057), .S(keyinput3), .Q(n974) );
  INVX0 U1315 ( .INP(n1252), .ZN(n1057) );
  NAND2X0 U1316 ( .IN1(N13), .IN2(N1), .QN(n1252) );
  NOR2X0 U1317 ( .IN1(n1081), .IN2(N13), .QN(n1286) );
  INVX0 U1318 ( .INP(N1), .ZN(n1081) );
  AO21X1 U1319 ( .IN1(n729), .IN2(n731), .IN3(n758), .Q(N1947) );
  INVX0 U1320 ( .INP(N87), .ZN(n758) );
  INVX0 U1321 ( .INP(N97), .ZN(n731) );
  INVX0 U1322 ( .INP(N107), .ZN(n729) );
endmodule

