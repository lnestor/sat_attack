`timescale 1ns / 1ps
// Verilog
// c432
// Ninputs 36
// Noutputs 7
// NtotalGates 160
// NOT1 40
// NAND2 64
// NOR2 19
// AND9 3
// XOR2 18
// NAND4 14
// AND8 1
// NAND3 1

module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
                  N430,N431,N432,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:56] KeyNOTWire_0;

input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;

output N223,N329,N370,N421,N430,N431,N432;

wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429;

  not NOT1_1 (KeyWire_0[0], N1);
  xor KeyGate_0_0(N118, keyIn_0_0, KeyWire_0[0]);
  not NOT1_2 (KeyWire_0[1], N4);
  xnor KeyGate_0_1(N119, keyIn_0_1, KeyWire_0[1]);
  not NOT1_3 (KeyWire_0[2], N11);
  xor KeyGate_0_2(N122, keyIn_0_2, KeyWire_0[2]);
  not NOT1_4 (KeyWire_0[3], N17);
  xor KeyGate_0_3(N123, keyIn_0_3, KeyWire_0[3]);
  not NOT1_5 (KeyWire_0[4], N24);
  xor KeyGate_0_4(KeyNOTWire_0[0], keyIn_0_4, KeyWire_0[4]);
  not KeyNOTGate_0_0(N126, KeyNOTWire_0[0]);
  not NOT1_6 (KeyWire_0[5], N30);
  xnor KeyGate_0_5(KeyNOTWire_0[1], keyIn_0_5, KeyWire_0[5]);
  not KeyNOTGate_0_1(N127, KeyNOTWire_0[1]);
  not NOT1_7 (KeyWire_0[6], N37);
  xnor KeyGate_0_6(N130, keyIn_0_6, KeyWire_0[6]);
not NOT1_8 (N131, N43);
  not NOT1_9 (KeyWire_0[7], N50);
  xor KeyGate_0_7(KeyNOTWire_0[2], keyIn_0_7, KeyWire_0[7]);
  not KeyNOTGate_0_2(N134, KeyNOTWire_0[2]);
  not NOT1_10 (KeyWire_0[8], N56);
  xor KeyGate_0_8(KeyNOTWire_0[3], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_3(N135, KeyNOTWire_0[3]);
not NOT1_11 (N138, N63);
not NOT1_12 (N139, N69);
  not NOT1_13 (KeyWire_0[9], N76);
  xnor KeyGate_0_9(KeyNOTWire_0[4], keyIn_0_9, KeyWire_0[9]);
  not KeyNOTGate_0_4(N142, KeyNOTWire_0[4]);
  not NOT1_14 (KeyWire_0[10], N82);
  xnor KeyGate_0_10(N143, keyIn_0_10, KeyWire_0[10]);
  not NOT1_15 (KeyWire_0[11], N89);
  xnor KeyGate_0_11(N146, keyIn_0_11, KeyWire_0[11]);
not NOT1_16 (N147, N95);
  not NOT1_17 (KeyWire_0[12], N102);
  xor KeyGate_0_12(KeyNOTWire_0[5], keyIn_0_12, KeyWire_0[12]);
  not KeyNOTGate_0_5(N150, KeyNOTWire_0[5]);
  not NOT1_18 (KeyWire_0[13], N108);
  xnor KeyGate_0_13(N151, keyIn_0_13, KeyWire_0[13]);
  nand NAND2_19 (KeyWire_0[14], N118, N4);
  xnor KeyGate_0_14(KeyNOTWire_0[6], keyIn_0_14, KeyWire_0[14]);
  not KeyNOTGate_0_6(N154, KeyNOTWire_0[6]);
  nor NOR2_20 (KeyWire_0[15], N8, N119);
  xor KeyGate_0_15(N157, keyIn_0_15, KeyWire_0[15]);
  nor NOR2_21 (KeyWire_0[16], N14, N119);
  xor KeyGate_0_16(N158, keyIn_0_16, KeyWire_0[16]);
nand NAND2_22 (N159, N122, N17);
  nand NAND2_23 (KeyWire_0[17], N126, N30);
  xor KeyGate_0_17(N162, keyIn_0_17, KeyWire_0[17]);
  nand NAND2_24 (KeyWire_0[18], N130, N43);
  xor KeyGate_0_18(N165, keyIn_0_18, KeyWire_0[18]);
  nand NAND2_25 (KeyWire_0[19], N134, N56);
  xor KeyGate_0_19(N168, keyIn_0_19, KeyWire_0[19]);
nand NAND2_26 (N171, N138, N69);
nand NAND2_27 (N174, N142, N82);
  nand NAND2_28 (KeyWire_0[20], N146, N95);
  xnor KeyGate_0_20(KeyNOTWire_0[7], keyIn_0_20, KeyWire_0[20]);
  not KeyNOTGate_0_7(N177, KeyNOTWire_0[7]);
  nand NAND2_29 (KeyWire_0[21], N150, N108);
  xnor KeyGate_0_21(KeyNOTWire_0[8], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_8(N180, KeyNOTWire_0[8]);
  nor NOR2_30 (KeyWire_0[22], N21, N123);
  xor KeyGate_0_22(N183, keyIn_0_22, KeyWire_0[22]);
nor NOR2_31 (N184, N27, N123);
  nor NOR2_32 (KeyWire_0[23], N34, N127);
  xnor KeyGate_0_23(KeyNOTWire_0[9], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_9(N185, KeyNOTWire_0[9]);
  nor NOR2_33 (KeyWire_0[24], N40, N127);
  xor KeyGate_0_24(N186, keyIn_0_24, KeyWire_0[24]);
  nor NOR2_34 (KeyWire_0[25], N47, N131);
  xor KeyGate_0_25(KeyNOTWire_0[10], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_10(N187, KeyNOTWire_0[10]);
  nor NOR2_35 (KeyWire_0[26], N53, N131);
  xnor KeyGate_0_26(KeyNOTWire_0[11], keyIn_0_26, KeyWire_0[26]);
  not KeyNOTGate_0_11(N188, KeyNOTWire_0[11]);
  nor NOR2_36 (KeyWire_0[27], N60, N135);
  xnor KeyGate_0_27(KeyNOTWire_0[12], keyIn_0_27, KeyWire_0[27]);
  not KeyNOTGate_0_12(N189, KeyNOTWire_0[12]);
  nor NOR2_37 (KeyWire_0[28], N66, N135);
  xnor KeyGate_0_28(N190, keyIn_0_28, KeyWire_0[28]);
  nor NOR2_38 (KeyWire_0[29], N73, N139);
  xor KeyGate_0_29(KeyNOTWire_0[13], keyIn_0_29, KeyWire_0[29]);
  not KeyNOTGate_0_13(N191, KeyNOTWire_0[13]);
  nor NOR2_39 (KeyWire_0[30], N79, N139);
  xnor KeyGate_0_30(N192, keyIn_0_30, KeyWire_0[30]);
  nor NOR2_40 (KeyWire_0[31], N86, N143);
  xor KeyGate_0_31(KeyNOTWire_0[14], keyIn_0_31, KeyWire_0[31]);
  not KeyNOTGate_0_14(N193, KeyNOTWire_0[14]);
  nor NOR2_41 (KeyWire_0[32], N92, N143);
  xnor KeyGate_0_32(N194, keyIn_0_32, KeyWire_0[32]);
  nor NOR2_42 (KeyWire_0[33], N99, N147);
  xor KeyGate_0_33(N195, keyIn_0_33, KeyWire_0[33]);
  nor NOR2_43 (KeyWire_0[34], N105, N147);
  xnor KeyGate_0_34(N196, keyIn_0_34, KeyWire_0[34]);
  nor NOR2_44 (KeyWire_0[35], N112, N151);
  xor KeyGate_0_35(KeyNOTWire_0[15], keyIn_0_35, KeyWire_0[35]);
  not KeyNOTGate_0_15(N197, KeyNOTWire_0[15]);
  nor NOR2_45 (KeyWire_0[36], N115, N151);
  xor KeyGate_0_36(N198, keyIn_0_36, KeyWire_0[36]);
and AND9_46 (N199, N154, N159, N162, N165, N168, N171, N174, N177, N180);
  not NOT1_47 (KeyWire_0[37], N199);
  xnor KeyGate_0_37(KeyNOTWire_0[16], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_16(N203, KeyNOTWire_0[16]);
not NOT1_48 (N213, N199);
  not NOT1_49 (KeyWire_0[38], N199);
  xnor KeyGate_0_38(N223, keyIn_0_38, KeyWire_0[38]);
xor XOR2_50 (N224, N203, N154);
  xor XOR2_51 (KeyWire_0[39], N203, N159);
  xor KeyGate_0_39(N227, keyIn_0_39, KeyWire_0[39]);
  xor XOR2_52 (KeyWire_0[40], N203, N162);
  xnor KeyGate_0_40(KeyNOTWire_0[17], keyIn_0_40, KeyWire_0[40]);
  not KeyNOTGate_0_17(N230, KeyNOTWire_0[17]);
  xor XOR2_53 (KeyWire_0[41], N203, N165);
  xnor KeyGate_0_41(KeyNOTWire_0[18], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_18(N233, KeyNOTWire_0[18]);
  xor XOR2_54 (KeyWire_0[42], N203, N168);
  xor KeyGate_0_42(KeyNOTWire_0[19], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_19(N236, KeyNOTWire_0[19]);
  xor XOR2_55 (KeyWire_0[43], N203, N171);
  xnor KeyGate_0_43(N239, keyIn_0_43, KeyWire_0[43]);
  nand NAND2_56 (KeyWire_0[44], N1, N213);
  xor KeyGate_0_44(KeyNOTWire_0[20], keyIn_0_44, KeyWire_0[44]);
  not KeyNOTGate_0_20(N242, KeyNOTWire_0[20]);
xor XOR2_57 (N243, N203, N174);
nand NAND2_58 (N246, N213, N11);
  xor XOR2_59 (KeyWire_0[45], N203, N177);
  xnor KeyGate_0_45(N247, keyIn_0_45, KeyWire_0[45]);
  nand NAND2_60 (KeyWire_0[46], N213, N24);
  xnor KeyGate_0_46(KeyNOTWire_0[21], keyIn_0_46, KeyWire_0[46]);
  not KeyNOTGate_0_21(N250, KeyNOTWire_0[21]);
  xor XOR2_61 (KeyWire_0[47], N203, N180);
  xor KeyGate_0_47(N251, keyIn_0_47, KeyWire_0[47]);
  nand NAND2_62 (KeyWire_0[48], N213, N37);
  xnor KeyGate_0_48(KeyNOTWire_0[22], keyIn_0_48, KeyWire_0[48]);
  not KeyNOTGate_0_22(N254, KeyNOTWire_0[22]);
  nand NAND2_63 (KeyWire_0[49], N213, N50);
  xor KeyGate_0_49(KeyNOTWire_0[23], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_23(N255, KeyNOTWire_0[23]);
  nand NAND2_64 (KeyWire_0[50], N213, N63);
  xnor KeyGate_0_50(N256, keyIn_0_50, KeyWire_0[50]);
  nand NAND2_65 (KeyWire_0[51], N213, N76);
  xnor KeyGate_0_51(N257, keyIn_0_51, KeyWire_0[51]);
  nand NAND2_66 (KeyWire_0[52], N213, N89);
  xor KeyGate_0_52(N258, keyIn_0_52, KeyWire_0[52]);
  nand NAND2_67 (KeyWire_0[53], N213, N102);
  xor KeyGate_0_53(N259, keyIn_0_53, KeyWire_0[53]);
  nand NAND2_68 (KeyWire_0[54], N224, N157);
  xnor KeyGate_0_54(KeyNOTWire_0[24], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_24(N260, KeyNOTWire_0[24]);
  nand NAND2_69 (KeyWire_0[55], N224, N158);
  xnor KeyGate_0_55(KeyNOTWire_0[25], keyIn_0_55, KeyWire_0[55]);
  not KeyNOTGate_0_25(N263, KeyNOTWire_0[25]);
  nand NAND2_70 (KeyWire_0[56], N227, N183);
  xnor KeyGate_0_56(N264, keyIn_0_56, KeyWire_0[56]);
  nand NAND2_71 (KeyWire_0[57], N230, N185);
  xor KeyGate_0_57(N267, keyIn_0_57, KeyWire_0[57]);
  nand NAND2_72 (KeyWire_0[58], N233, N187);
  xor KeyGate_0_58(KeyNOTWire_0[26], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_26(N270, KeyNOTWire_0[26]);
nand NAND2_73 (N273, N236, N189);
  nand NAND2_74 (KeyWire_0[59], N239, N191);
  xor KeyGate_0_59(N276, keyIn_0_59, KeyWire_0[59]);
  nand NAND2_75 (KeyWire_0[60], N243, N193);
  xor KeyGate_0_60(KeyNOTWire_0[27], keyIn_0_60, KeyWire_0[60]);
  not KeyNOTGate_0_27(N279, KeyNOTWire_0[27]);
  nand NAND2_76 (KeyWire_0[61], N247, N195);
  xor KeyGate_0_61(N282, keyIn_0_61, KeyWire_0[61]);
  nand NAND2_77 (KeyWire_0[62], N251, N197);
  xnor KeyGate_0_62(N285, keyIn_0_62, KeyWire_0[62]);
  nand NAND2_78 (KeyWire_0[63], N227, N184);
  xor KeyGate_0_63(KeyNOTWire_0[28], keyIn_0_63, KeyWire_0[63]);
  not KeyNOTGate_0_28(N288, KeyNOTWire_0[28]);
  nand NAND2_79 (KeyWire_0[64], N230, N186);
  xnor KeyGate_0_64(KeyNOTWire_0[29], keyIn_0_64, KeyWire_0[64]);
  not KeyNOTGate_0_29(N289, KeyNOTWire_0[29]);
  nand NAND2_80 (KeyWire_0[65], N233, N188);
  xor KeyGate_0_65(N290, keyIn_0_65, KeyWire_0[65]);
  nand NAND2_81 (KeyWire_0[66], N236, N190);
  xor KeyGate_0_66(KeyNOTWire_0[30], keyIn_0_66, KeyWire_0[66]);
  not KeyNOTGate_0_30(N291, KeyNOTWire_0[30]);
  nand NAND2_82 (KeyWire_0[67], N239, N192);
  xor KeyGate_0_67(N292, keyIn_0_67, KeyWire_0[67]);
  nand NAND2_83 (KeyWire_0[68], N243, N194);
  xor KeyGate_0_68(KeyNOTWire_0[31], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_31(N293, KeyNOTWire_0[31]);
  nand NAND2_84 (KeyWire_0[69], N247, N196);
  xnor KeyGate_0_69(N294, keyIn_0_69, KeyWire_0[69]);
  nand NAND2_85 (KeyWire_0[70], N251, N198);
  xor KeyGate_0_70(KeyNOTWire_0[32], keyIn_0_70, KeyWire_0[70]);
  not KeyNOTGate_0_32(N295, KeyNOTWire_0[32]);
  and AND9_86 (KeyWire_0[71], N260, N264, N267, N270, N273, N276, N279, N282, N285);
  xnor KeyGate_0_71(N296, keyIn_0_71, KeyWire_0[71]);
  not NOT1_87 (KeyWire_0[72], N263);
  xor KeyGate_0_72(KeyNOTWire_0[33], keyIn_0_72, KeyWire_0[72]);
  not KeyNOTGate_0_33(N300, KeyNOTWire_0[33]);
not NOT1_88 (N301, N288);
  not NOT1_89 (KeyWire_0[73], N289);
  xnor KeyGate_0_73(N302, keyIn_0_73, KeyWire_0[73]);
not NOT1_90 (N303, N290);
not NOT1_91 (N304, N291);
  not NOT1_92 (KeyWire_0[74], N292);
  xor KeyGate_0_74(N305, keyIn_0_74, KeyWire_0[74]);
  not NOT1_93 (KeyWire_0[75], N293);
  xor KeyGate_0_75(N306, keyIn_0_75, KeyWire_0[75]);
  not NOT1_94 (KeyWire_0[76], N294);
  xnor KeyGate_0_76(KeyNOTWire_0[34], keyIn_0_76, KeyWire_0[76]);
  not KeyNOTGate_0_34(N307, KeyNOTWire_0[34]);
  not NOT1_95 (KeyWire_0[77], N295);
  xnor KeyGate_0_77(N308, keyIn_0_77, KeyWire_0[77]);
  not NOT1_96 (KeyWire_0[78], N296);
  xor KeyGate_0_78(KeyNOTWire_0[35], keyIn_0_78, KeyWire_0[78]);
  not KeyNOTGate_0_35(N309, KeyNOTWire_0[35]);
  not NOT1_97 (KeyWire_0[79], N296);
  xnor KeyGate_0_79(KeyNOTWire_0[36], keyIn_0_79, KeyWire_0[79]);
  not KeyNOTGate_0_36(N319, KeyNOTWire_0[36]);
  not NOT1_98 (KeyWire_0[80], N296);
  xnor KeyGate_0_80(N329, keyIn_0_80, KeyWire_0[80]);
  xor XOR2_99 (KeyWire_0[81], N309, N260);
  xor KeyGate_0_81(KeyNOTWire_0[37], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_37(N330, KeyNOTWire_0[37]);
  xor XOR2_100 (KeyWire_0[82], N309, N264);
  xor KeyGate_0_82(KeyNOTWire_0[38], keyIn_0_82, KeyWire_0[82]);
  not KeyNOTGate_0_38(N331, KeyNOTWire_0[38]);
xor XOR2_101 (N332, N309, N267);
xor XOR2_102 (N333, N309, N270);
nand NAND2_103 (N334, N8, N319);
  xor XOR2_104 (KeyWire_0[83], N309, N273);
  xor KeyGate_0_83(N335, keyIn_0_83, KeyWire_0[83]);
  nand NAND2_105 (KeyWire_0[84], N319, N21);
  xnor KeyGate_0_84(KeyNOTWire_0[39], keyIn_0_84, KeyWire_0[84]);
  not KeyNOTGate_0_39(N336, KeyNOTWire_0[39]);
  xor XOR2_106 (KeyWire_0[85], N309, N276);
  xor KeyGate_0_85(KeyNOTWire_0[40], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_40(N337, KeyNOTWire_0[40]);
nand NAND2_107 (N338, N319, N34);
  xor XOR2_108 (KeyWire_0[86], N309, N279);
  xnor KeyGate_0_86(N339, keyIn_0_86, KeyWire_0[86]);
  nand NAND2_109 (KeyWire_0[87], N319, N47);
  xor KeyGate_0_87(KeyNOTWire_0[41], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_41(N340, KeyNOTWire_0[41]);
  xor XOR2_110 (KeyWire_0[88], N309, N282);
  xnor KeyGate_0_88(N341, keyIn_0_88, KeyWire_0[88]);
  nand NAND2_111 (KeyWire_0[89], N319, N60);
  xnor KeyGate_0_89(N342, keyIn_0_89, KeyWire_0[89]);
  xor XOR2_112 (KeyWire_0[90], N309, N285);
  xor KeyGate_0_90(N343, keyIn_0_90, KeyWire_0[90]);
  nand NAND2_113 (KeyWire_0[91], N319, N73);
  xnor KeyGate_0_91(N344, keyIn_0_91, KeyWire_0[91]);
nand NAND2_114 (N345, N319, N86);
  nand NAND2_115 (KeyWire_0[92], N319, N99);
  xor KeyGate_0_92(KeyNOTWire_0[42], keyIn_0_92, KeyWire_0[92]);
  not KeyNOTGate_0_42(N346, KeyNOTWire_0[42]);
nand NAND2_116 (N347, N319, N112);
  nand NAND2_117 (KeyWire_0[93], N330, N300);
  xor KeyGate_0_93(N348, keyIn_0_93, KeyWire_0[93]);
  nand NAND2_118 (KeyWire_0[94], N331, N301);
  xor KeyGate_0_94(KeyNOTWire_0[43], keyIn_0_94, KeyWire_0[94]);
  not KeyNOTGate_0_43(N349, KeyNOTWire_0[43]);
  nand NAND2_119 (KeyWire_0[95], N332, N302);
  xor KeyGate_0_95(N350, keyIn_0_95, KeyWire_0[95]);
  nand NAND2_120 (KeyWire_0[96], N333, N303);
  xnor KeyGate_0_96(N351, keyIn_0_96, KeyWire_0[96]);
nand NAND2_121 (N352, N335, N304);
  nand NAND2_122 (KeyWire_0[97], N337, N305);
  xnor KeyGate_0_97(N353, keyIn_0_97, KeyWire_0[97]);
nand NAND2_123 (N354, N339, N306);
  nand NAND2_124 (KeyWire_0[98], N341, N307);
  xor KeyGate_0_98(N355, keyIn_0_98, KeyWire_0[98]);
  nand NAND2_125 (KeyWire_0[99], N343, N308);
  xnor KeyGate_0_99(N356, keyIn_0_99, KeyWire_0[99]);
and AND9_126 (N357, N348, N349, N350, N351, N352, N353, N354, N355, N356);
  not NOT1_127 (KeyWire_0[100], N357);
  xnor KeyGate_0_100(KeyNOTWire_0[44], keyIn_0_100, KeyWire_0[100]);
  not KeyNOTGate_0_44(N360, KeyNOTWire_0[44]);
not NOT1_128 (N370, N357);
  nand NAND2_129 (KeyWire_0[101], N14, N360);
  xor KeyGate_0_101(KeyNOTWire_0[45], keyIn_0_101, KeyWire_0[101]);
  not KeyNOTGate_0_45(N371, KeyNOTWire_0[45]);
  nand NAND2_130 (KeyWire_0[102], N360, N27);
  xnor KeyGate_0_102(N372, keyIn_0_102, KeyWire_0[102]);
  nand NAND2_131 (KeyWire_0[103], N360, N40);
  xnor KeyGate_0_103(N373, keyIn_0_103, KeyWire_0[103]);
  nand NAND2_132 (KeyWire_0[104], N360, N53);
  xor KeyGate_0_104(N374, keyIn_0_104, KeyWire_0[104]);
  nand NAND2_133 (KeyWire_0[105], N360, N66);
  xnor KeyGate_0_105(KeyNOTWire_0[46], keyIn_0_105, KeyWire_0[105]);
  not KeyNOTGate_0_46(N375, KeyNOTWire_0[46]);
  nand NAND2_134 (KeyWire_0[106], N360, N79);
  xor KeyGate_0_106(N376, keyIn_0_106, KeyWire_0[106]);
  nand NAND2_135 (KeyWire_0[107], N360, N92);
  xnor KeyGate_0_107(N377, keyIn_0_107, KeyWire_0[107]);
  nand NAND2_136 (KeyWire_0[108], N360, N105);
  xor KeyGate_0_108(N378, keyIn_0_108, KeyWire_0[108]);
nand NAND2_137 (N379, N360, N115);
  nand NAND4_138 (KeyWire_0[109], N4, N242, N334, N371);
  xor KeyGate_0_109(KeyNOTWire_0[47], keyIn_0_109, KeyWire_0[109]);
  not KeyNOTGate_0_47(N380, KeyNOTWire_0[47]);
  nand NAND4_139 (KeyWire_0[110], N246, N336, N372, N17);
  xnor KeyGate_0_110(N381, keyIn_0_110, KeyWire_0[110]);
  nand NAND4_140 (KeyWire_0[111], N250, N338, N373, N30);
  xnor KeyGate_0_111(KeyNOTWire_0[48], keyIn_0_111, KeyWire_0[111]);
  not KeyNOTGate_0_48(N386, KeyNOTWire_0[48]);
nand NAND4_141 (N393, N254, N340, N374, N43);
  nand NAND4_142 (KeyWire_0[112], N255, N342, N375, N56);
  xnor KeyGate_0_112(N399, keyIn_0_112, KeyWire_0[112]);
  nand NAND4_143 (KeyWire_0[113], N256, N344, N376, N69);
  xnor KeyGate_0_113(KeyNOTWire_0[49], keyIn_0_113, KeyWire_0[113]);
  not KeyNOTGate_0_49(N404, KeyNOTWire_0[49]);
  nand NAND4_144 (KeyWire_0[114], N257, N345, N377, N82);
  xor KeyGate_0_114(N407, keyIn_0_114, KeyWire_0[114]);
nand NAND4_145 (N411, N258, N346, N378, N95);
nand NAND4_146 (N414, N259, N347, N379, N108);
not NOT1_147 (N415, N380);
  and AND8_148 (KeyWire_0[115], N381, N386, N393, N399, N404, N407, N411, N414);
  xor KeyGate_0_115(KeyNOTWire_0[50], keyIn_0_115, KeyWire_0[115]);
  not KeyNOTGate_0_50(N416, KeyNOTWire_0[50]);
  not NOT1_149 (KeyWire_0[116], N393);
  xor KeyGate_0_116(KeyNOTWire_0[51], keyIn_0_116, KeyWire_0[116]);
  not KeyNOTGate_0_51(N417, KeyNOTWire_0[51]);
  not NOT1_150 (KeyWire_0[117], N404);
  xor KeyGate_0_117(N418, keyIn_0_117, KeyWire_0[117]);
  not NOT1_151 (KeyWire_0[118], N407);
  xnor KeyGate_0_118(KeyNOTWire_0[52], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_52(N419, KeyNOTWire_0[52]);
  not NOT1_152 (KeyWire_0[119], N411);
  xor KeyGate_0_119(KeyNOTWire_0[53], keyIn_0_119, KeyWire_0[119]);
  not KeyNOTGate_0_53(N420, KeyNOTWire_0[53]);
  nor NOR2_153 (KeyWire_0[120], N415, N416);
  xnor KeyGate_0_120(KeyNOTWire_0[54], keyIn_0_120, KeyWire_0[120]);
  not KeyNOTGate_0_54(N421, KeyNOTWire_0[54]);
  nand NAND2_154 (KeyWire_0[121], N386, N417);
  xor KeyGate_0_121(KeyNOTWire_0[55], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_55(N422, KeyNOTWire_0[55]);
  nand NAND4_155 (KeyWire_0[122], N386, N393, N418, N399);
  xnor KeyGate_0_122(KeyNOTWire_0[56], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_56(N425, KeyNOTWire_0[56]);
  nand NAND3_156 (KeyWire_0[123], N399, N393, N419);
  xor KeyGate_0_123(N428, keyIn_0_123, KeyWire_0[123]);
  nand NAND4_157 (KeyWire_0[124], N386, N393, N407, N420);
  xor KeyGate_0_124(N429, keyIn_0_124, KeyWire_0[124]);
  nand NAND4_158 (KeyWire_0[125], N381, N386, N422, N399);
  xor KeyGate_0_125(N430, keyIn_0_125, KeyWire_0[125]);
  nand NAND4_159 (KeyWire_0[126], N381, N386, N425, N428);
  xnor KeyGate_0_126(N431, keyIn_0_126, KeyWire_0[126]);
  nand NAND4_160 (KeyWire_0[127], N381, N422, N425, N429);
  xnor KeyGate_0_127(N432, keyIn_0_127, KeyWire_0[127]);

endmodule
