
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47,
         N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92,
         N95, N99, N102, N105, N108, N112, N115, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284;

  XNOR2X1 U151 ( .IN1(keyinput31), .IN2(n149), .Q(N432) );
  OA21X1 U152 ( .IN1(n150), .IN2(n151), .IN3(n152), .Q(n149) );
  OA221X1 U153 ( .IN1(n153), .IN2(n154), .IN3(n155), .IN4(n156), .IN5(n157), 
        .Q(n150) );
  INVX0 U154 ( .INP(n158), .ZN(n155) );
  INVX0 U155 ( .INP(n159), .ZN(n153) );
  NAND3X0 U156 ( .IN1(n160), .IN2(n152), .IN3(n161), .QN(N431) );
  NAND3X0 U157 ( .IN1(n157), .IN2(n158), .IN3(n162), .QN(n160) );
  XNOR2X1 U158 ( .IN1(keyinput30), .IN2(n163), .Q(N430) );
  NOR2X0 U159 ( .IN1(n164), .IN2(n165), .QN(N421) );
  OA221X1 U160 ( .IN1(n166), .IN2(n167), .IN3(n168), .IN4(n169), .IN5(n170), 
        .Q(n165) );
  OA21X1 U161 ( .IN1(n171), .IN2(n172), .IN3(N4), .Q(n170) );
  INVX0 U162 ( .INP(N1), .ZN(n169) );
  NOR4X0 U163 ( .IN1(n173), .IN2(n174), .IN3(n163), .IN4(n162), .QN(n164) );
  NAND2X0 U164 ( .IN1(n156), .IN2(n159), .QN(n162) );
  AO221X1 U165 ( .IN1(N86), .IN2(N329), .IN3(N92), .IN4(N370), .IN5(n175), .Q(
        n159) );
  MUX21X1 U166 ( .IN1(n176), .IN2(n177), .S(keyinput15), .Q(n175) );
  NAND3X0 U167 ( .IN1(N76), .IN2(N82), .IN3(n178), .QN(n177) );
  AO21X1 U168 ( .IN1(n178), .IN2(N76), .IN3(n179), .Q(n176) );
  XOR2X1 U169 ( .IN1(n180), .IN2(keyinput29), .Q(n156) );
  NAND3X0 U170 ( .IN1(n181), .IN2(n182), .IN3(n183), .QN(n180) );
  XOR2X1 U171 ( .IN1(n184), .IN2(keyinput27), .Q(n183) );
  NAND2X0 U172 ( .IN1(N79), .IN2(N370), .QN(n184) );
  AO21X1 U173 ( .IN1(N69), .IN2(n168), .IN3(n185), .Q(n182) );
  XOR2X1 U174 ( .IN1(n186), .IN2(keyinput24), .Q(n181) );
  NAND4X0 U175 ( .IN1(n161), .IN2(n157), .IN3(n158), .IN4(n152), .QN(n163) );
  AO222X1 U176 ( .IN1(N21), .IN2(N329), .IN3(n187), .IN4(n188), .IN5(N27), 
        .IN6(N370), .Q(n152) );
  NAND2X0 U177 ( .IN1(N17), .IN2(n168), .QN(n187) );
  AO221X1 U178 ( .IN1(n178), .IN2(N50), .IN3(N60), .IN4(N329), .IN5(n189), .Q(
        n158) );
  AO21X1 U179 ( .IN1(N66), .IN2(N370), .IN3(n190), .Q(n189) );
  INVX0 U180 ( .INP(n168), .ZN(n178) );
  AO222X1 U181 ( .IN1(N47), .IN2(N329), .IN3(n191), .IN4(n192), .IN5(N53), 
        .IN6(N370), .Q(n157) );
  NAND2X0 U182 ( .IN1(N43), .IN2(n168), .QN(n191) );
  INVX0 U183 ( .INP(n151), .ZN(n161) );
  XNOR2X1 U184 ( .IN1(n193), .IN2(keyinput28), .Q(n151) );
  AO222X1 U185 ( .IN1(N34), .IN2(N329), .IN3(n194), .IN4(n195), .IN5(N40), 
        .IN6(N370), .Q(n193) );
  NAND2X0 U186 ( .IN1(N30), .IN2(n168), .QN(n194) );
  INVX0 U187 ( .INP(n154), .ZN(n174) );
  AO221X1 U188 ( .IN1(n196), .IN2(n197), .IN3(N105), .IN4(N370), .IN5(n198), 
        .Q(n154) );
  XOR2X1 U189 ( .IN1(keyinput25), .IN2(n199), .Q(n198) );
  NOR2X0 U190 ( .IN1(n166), .IN2(n200), .QN(n199) );
  NAND2X0 U191 ( .IN1(N95), .IN2(n168), .QN(n196) );
  OA221X1 U192 ( .IN1(n166), .IN2(n201), .IN3(n171), .IN4(n202), .IN5(n203), 
        .Q(n173) );
  OA21X1 U193 ( .IN1(n168), .IN2(n204), .IN3(N108), .Q(n203) );
  XNOR2X1 U194 ( .IN1(N223), .IN2(keyinput9), .Q(n168) );
  INVX0 U195 ( .INP(N370), .ZN(n171) );
  NAND4X0 U196 ( .IN1(n205), .IN2(n206), .IN3(n207), .IN4(n208), .QN(N370) );
  NOR4X0 U197 ( .IN1(n209), .IN2(n210), .IN3(n211), .IN4(n212), .QN(n208) );
  XOR2X1 U198 ( .IN1(n213), .IN2(keyinput26), .Q(n212) );
  OR3X1 U199 ( .IN1(n214), .IN2(N27), .IN3(n215), .Q(n213) );
  NOR2X0 U200 ( .IN1(n166), .IN2(n216), .QN(n214) );
  NOR2X0 U201 ( .IN1(n217), .IN2(n218), .QN(n211) );
  XOR2X1 U202 ( .IN1(n219), .IN2(keyinput20), .Q(n218) );
  NAND2X0 U203 ( .IN1(n220), .IN2(n221), .QN(n219) );
  XOR2X1 U204 ( .IN1(keyinput5), .IN2(n222), .Q(n220) );
  NOR2X0 U205 ( .IN1(N40), .IN2(n223), .QN(n222) );
  XNOR3X1 U206 ( .IN1(keyinput23), .IN2(n224), .IN3(N329), .Q(n217) );
  OA21X1 U207 ( .IN1(n166), .IN2(n225), .IN3(n226), .Q(n210) );
  XOR2X1 U208 ( .IN1(n227), .IN2(keyinput19), .Q(n226) );
  NAND2X0 U209 ( .IN1(n228), .IN2(n202), .QN(n227) );
  INVX0 U210 ( .INP(N115), .ZN(n202) );
  OA21X1 U211 ( .IN1(n229), .IN2(n166), .IN3(n230), .Q(n209) );
  XOR2X1 U212 ( .IN1(n231), .IN2(keyinput21), .Q(n230) );
  OR2X1 U213 ( .IN1(n232), .IN2(N66), .Q(n231) );
  AND3X1 U214 ( .IN1(n233), .IN2(n234), .IN3(n235), .Q(n207) );
  NAND4X0 U215 ( .IN1(N69), .IN2(n236), .IN3(n186), .IN4(n237), .QN(n235) );
  INVX0 U216 ( .INP(N79), .ZN(n237) );
  NAND2X0 U217 ( .IN1(N73), .IN2(N329), .QN(n186) );
  OR3X1 U218 ( .IN1(n238), .IN2(N92), .IN3(n239), .Q(n234) );
  NOR2X0 U219 ( .IN1(n166), .IN2(n240), .QN(n238) );
  NAND4X0 U220 ( .IN1(n241), .IN2(n242), .IN3(n243), .IN4(n172), .QN(n233) );
  INVX0 U221 ( .INP(N14), .ZN(n172) );
  XNOR3X1 U222 ( .IN1(keyinput22), .IN2(n244), .IN3(N329), .Q(n241) );
  NAND3X0 U223 ( .IN1(n245), .IN2(n246), .IN3(n247), .QN(n206) );
  XOR2X1 U224 ( .IN1(n248), .IN2(keyinput8), .Q(n247) );
  NAND2X0 U225 ( .IN1(n249), .IN2(n250), .QN(n248) );
  INVX0 U226 ( .INP(N105), .ZN(n250) );
  NAND2X0 U227 ( .IN1(n251), .IN2(N329), .QN(n245) );
  NAND3X0 U228 ( .IN1(n252), .IN2(n253), .IN3(n254), .QN(n205) );
  XOR2X1 U229 ( .IN1(n255), .IN2(keyinput7), .Q(n254) );
  OR2X1 U230 ( .IN1(n256), .IN2(N53), .Q(n255) );
  NAND2X0 U231 ( .IN1(N329), .IN2(n257), .QN(n253) );
  INVX0 U232 ( .INP(n166), .ZN(N329) );
  NOR4X0 U233 ( .IN1(n216), .IN2(n240), .IN3(n258), .IN4(n259), .QN(n166) );
  NAND4X0 U234 ( .IN1(n224), .IN2(n251), .IN3(n260), .IN4(n261), .QN(n259) );
  NAND3X0 U235 ( .IN1(n236), .IN2(n262), .IN3(N69), .QN(n261) );
  INVX0 U236 ( .INP(N73), .ZN(n262) );
  XNOR3X1 U237 ( .IN1(keyinput13), .IN2(n185), .IN3(N223), .Q(n236) );
  INVX0 U238 ( .INP(n225), .ZN(n260) );
  XNOR2X1 U239 ( .IN1(n263), .IN2(keyinput18), .Q(n225) );
  NAND2X0 U240 ( .IN1(n228), .IN2(n201), .QN(n263) );
  INVX0 U241 ( .INP(N112), .ZN(n201) );
  AND2X1 U242 ( .IN1(n264), .IN2(n265), .Q(n228) );
  XOR3X1 U243 ( .IN1(keyinput14), .IN2(n266), .IN3(N223), .Q(n265) );
  XNOR2X1 U244 ( .IN1(N108), .IN2(keyinput3), .Q(n264) );
  XOR2X1 U245 ( .IN1(n267), .IN2(keyinput17), .Q(n251) );
  NAND3X0 U246 ( .IN1(n246), .IN2(n200), .IN3(n249), .QN(n267) );
  XOR2X1 U247 ( .IN1(N95), .IN2(keyinput2), .Q(n249) );
  INVX0 U248 ( .INP(N99), .ZN(n200) );
  NAND2X0 U249 ( .IN1(N223), .IN2(n197), .QN(n246) );
  XOR2X1 U250 ( .IN1(n268), .IN2(keyinput16), .Q(n224) );
  NAND3X0 U251 ( .IN1(n221), .IN2(n269), .IN3(N30), .QN(n268) );
  INVX0 U252 ( .INP(N34), .ZN(n269) );
  XOR3X1 U253 ( .IN1(keyinput11), .IN2(n195), .IN3(N223), .Q(n221) );
  NAND3X0 U254 ( .IN1(n257), .IN2(n270), .IN3(n244), .QN(n258) );
  NAND3X0 U255 ( .IN1(n243), .IN2(n167), .IN3(n242), .QN(n244) );
  XNOR2X1 U256 ( .IN1(n271), .IN2(keyinput0), .Q(n242) );
  INVX0 U257 ( .INP(N8), .ZN(n167) );
  OAI21X1 U258 ( .IN1(n271), .IN2(N1), .IN3(N223), .QN(n243) );
  INVX0 U259 ( .INP(n229), .ZN(n270) );
  NOR2X0 U260 ( .IN1(n232), .IN2(N60), .QN(n229) );
  AO21X1 U261 ( .IN1(N50), .IN2(N223), .IN3(n190), .Q(n232) );
  NAND2X0 U262 ( .IN1(n272), .IN2(n252), .QN(n257) );
  XNOR3X1 U263 ( .IN1(keyinput12), .IN2(n192), .IN3(N223), .Q(n252) );
  INVX0 U264 ( .INP(n273), .ZN(n192) );
  XOR2X1 U265 ( .IN1(n274), .IN2(keyinput6), .Q(n272) );
  OR2X1 U266 ( .IN1(n256), .IN2(N47), .Q(n274) );
  NOR2X0 U267 ( .IN1(n239), .IN2(N86), .QN(n240) );
  AO21X1 U268 ( .IN1(N76), .IN2(N223), .IN3(n179), .Q(n239) );
  NOR2X0 U269 ( .IN1(n215), .IN2(N21), .QN(n216) );
  NAND2X0 U270 ( .IN1(n275), .IN2(n276), .QN(n215) );
  XNOR3X1 U271 ( .IN1(keyinput10), .IN2(n188), .IN3(N223), .Q(n276) );
  INVX0 U272 ( .INP(n277), .ZN(n188) );
  XOR2X1 U273 ( .IN1(n278), .IN2(keyinput1), .Q(n275) );
  NAND4X0 U274 ( .IN1(n197), .IN2(n195), .IN3(n279), .IN4(n280), .QN(N223) );
  OA221X1 U275 ( .IN1(N50), .IN2(n190), .IN3(N1), .IN4(n271), .IN5(n281), .Q(
        n280) );
  OA21X1 U276 ( .IN1(N76), .IN2(n179), .IN3(n266), .Q(n281) );
  XNOR2X1 U277 ( .IN1(n282), .IN2(keyinput4), .Q(n266) );
  NAND2X0 U278 ( .IN1(N108), .IN2(n204), .QN(n282) );
  INVX0 U279 ( .INP(N102), .ZN(n204) );
  INVX0 U280 ( .INP(N82), .ZN(n179) );
  INVX0 U281 ( .INP(N4), .ZN(n271) );
  INVX0 U282 ( .INP(N56), .ZN(n190) );
  NOR3X0 U283 ( .IN1(n277), .IN2(n185), .IN3(n273), .QN(n279) );
  NOR2X0 U284 ( .IN1(N37), .IN2(n256), .QN(n273) );
  INVX0 U285 ( .INP(N43), .ZN(n256) );
  NOR2X0 U286 ( .IN1(N63), .IN2(n283), .QN(n185) );
  INVX0 U287 ( .INP(N69), .ZN(n283) );
  NOR2X0 U288 ( .IN1(N11), .IN2(n278), .QN(n277) );
  INVX0 U289 ( .INP(N17), .ZN(n278) );
  OR2X1 U290 ( .IN1(N24), .IN2(n223), .Q(n195) );
  INVX0 U291 ( .INP(N30), .ZN(n223) );
  NAND2X0 U292 ( .IN1(n284), .IN2(N95), .QN(n197) );
  INVX0 U293 ( .INP(N89), .ZN(n284) );
endmodule

