// Verilog File 
module c1908.bench (G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953,G3,G6,G9,G12,G30,G45,
G48,G15,G18,G21,G24,G27,G33,G36,G39,G42,
G75,G51,G54,G60,G63,G66,G69,G72,G57);

input G101,G104,G107,G110,G113,G116,G119,G122,G125,
G128,G131,G134,G137,G140,G143,G146,G210,G214,G217,
G221,G224,G227,G234,G237,G469,G472,G475,G478,G898,
G900,G902,G952,G953;


output G3, G6, G9, G12, G30, G45, G48, G15, G18, 
G21, G24, G27, G33, G36, G39, G42, G75, G51, G54, 
G60, G63, G66, G69, G72, G57;

wire G149, G153, G156, G160, G165, G168, G171, G175, G179, 
G184, G188, G191, G194, G198, G202, G206, G231, G233, G241, 
G244, G245, G248, G517, G529, G541, G553, G859, G862, G907, 
G909, G911, G918, G919, G922, G926, G930, G932, G934, G938, 
G943, G947, G949, G1506, G1514, G1522, G1530, G1538, G1546, G1554, 
G1562, G1570, G1578, G1586, G1594, G1602, G1610, G1618, G1626, G1512, 
G1520, G1528, G1536, G1544, G1552, G1560, G1568, G1576, G1584, G1592, 
G1600, G1608, G1616, G1624, G1632, G50, G52, G56, G58, G62, 
G64, G251, G254, G288, G291, G299, G302, G318, G321, G327, 
G330, G352, G355, G369, G382, G385, G853, G856, G893, G954, 
G955, G1050, G1053, G1176, G1179, G1197, G1207, G1222, G1244, G1278, 
G1290, G1300, G1312, G1332, G1335, G1442, G1450, G1458, G1466, G1474, 
G1482, G1490, G1498, G1634, G1644, G1657, G1665, G1697, G1705, G1713, 
G1721, G1745, G1753, G1785, G1793, G1814, G1817, G1830, G1833, G1841, 
G1849, G1854, G1857, G1870, G1873, G1878, G1881, G1642, G1652, G1056, 
G1057, G1182, G1183, G1211, G1298, G1320, G1338, G1339, G457, G459, 
G482, G487, G492, G505, G1456, G1448, G1472, G1464, G1488, G1480, 
G1504, G1496, G956, G967, G978, G979, G980, G1661, G990, G1669, 
G1030, G1701, G1040, G1709, G1058, G1717, G1068, G1725, G1078, G1090, 
G1100, G1749, G1112, G1757, G1154, G1789, G1166, G1797, G1194, G1201, 
G1204, G1820, G1821, G1230, G1836, G1837, G1252, G1256, G1845, G1268, 
G1853, G1860, G1861, G1286, G1876, G1877, G1308, G1884, G1885, G1654, 
G1662, G1694, G1702, G1710, G1718, G1726, G1734, G1742, G1750, G1782, 
G1790, G1838, G1846, G297, G298, G361, G362, G404, G405, G1225, 
G1226, G1247, G1248, G1281, G1282, G1303, G1304, G1315, G1316, G998, 
G988, G268, G1038, G1048, G1076, G1066, G1098, G1120, G1174, G363, 
G1210, G373, G1276, G406, G565, G566, G614, G615, G958, G969, 
G1660, G984, G1668, G994, G1700, G1034, G1708, G1044, G1716, G1062, 
G1724, G1072, G1732, G1086, G1740, G1748, G1104, G1108, G1756, G1116, 
G1788, G1158, G1162, G1796, G1170, G1200, G1203, G1227, G1249, G1844, 
G1260, G1264, G1852, G1272, G1283, G1305, G1317, G1410, G1418, G1426, 
G1434, G269, G372, G983, G993, G1033, G1043, G1061, G1071, G1103, 
G1115, G1157, G1169, G1184, G1202, G1259, G1271, G1322, G374, G396, 
G1321, G1424, G1416, G1440, G1432, G985, G995, G1035, G1045, G1063, 
G1073, G1105, G1117, G1159, G1171, G1212, G1231, G1232, G1253, G1254, 
G1261, G1273, G1287, G1288, G1309, G1310, G1192, G397, G1330, G1000, 
G1010, G1233, G1255, G1289, G1311, G1381, G257, G999, G260, G989, 
G272, G1039, G294, G1049, G305, G1077, G308, G1067, G333, G1121, 
G358, G1175, G1220, G388, G1277, G398, G1109, G1110, G1163, G1164, 
G1234, G1265, G1266, G1822, G1862, G1865, G258, G261, G273, G1018, 
G1008, G295, G306, G309, G334, G359, G389, G1385, G1111, G1165, 
G1267, G1886, G259, G262, G274, G296, G307, G310, G335, G360, 
G1242, G390, G1828, G1868, G1869, G1373, G1798, G1825, G265, G314, 
G336, G407, G1293, G1294, G1892, G1777, G1889, G410, G1377, G1804, 
G1237, G1829, G1295, G1670, G1678, G1729, G1737, G1761, G1769, G340, 
G343, G1781, G1238, G1325, G1893, G1340, G1352, G1673, G1681, G1801, 
G1897, G1905, G391, G1299, G1676, G1684, G1081, G1733, G1093, G1741, 
G1765, G1773, G1239, G1326, G1894, G1902, G392, G1360, G1003, G1677, 
G1013, G1685, G1082, G1094, G1122, G1134, G1187, G1805, G1327, G1901, 
G1348, G1909, G1758, G1766, G377, G1243, G393, G1004, G1014, G1083, 
G1095, G1188, G1900, G1344, G1908, G1356, G1142, G378, G399, G1331, 
G1005, G1015, G1764, G1126, G1130, G1772, G1138, G1189, G1343, G1355, 
G324, G1099, G379, G400, G449, G1087, G1088, G1125, G1137, G1345, 
G1357, G1397, G277, G1019, G280, G1009, G325, G364, G1193, G401, 
G1089, G1127, G1139, G278, G281, G326, G365, G413, G1361, G1401, 
G445, G1349, G1350, G1389, G1493, G1501, G1689, G279, G282, G346, 
G1143, G366, G414, G453, G1131, G1132, G1351, G1365, G1405, G285, 
G347, G367, G415, G1393, G556, G1505, G559, G1497, G1693, G1133, 
G1477, G1485, G1809, G348, G1369, G1409, G557, G560, G1362, G1378, 
G1429, G1437, G1686, G1774, G1910, G1918, G544, G1489, G547, G1481, 
G558, G561, G1813, G1370, G1368, G417, G1384, G424, G508, G1441, 
G511, G1433, G545, G548, G564, G1692, G1024, G1780, G1148, G1916, 
G1924, G416, G1376, G421, G423, G509, G512, G546, G549, G719, 
G722, G1023, G1147, G418, G420, G425, G510, G513, G552, G1025, 
G1149, G419, G422, G441, G516, G725, G728, G1029, G1153, G433, 
G437, G663, G666, G731, G746, G756, G770, G1461, G1469, G1413, 
G1421, G1445, G1453, G532, G1473, G535, G1465, G495, G1425, G498, 
G1417, G520, G1457, G523, G1449, G533, G536, G496, G499, G521, 
G524, G534, G537, G497, G500, G522, G525, G540, G503, G528, 
G669, G672, G569, G588, G618, G639, G867, G588a, G588b, G639a, 
G639b, G675, G688, G696, G710, G73, G572, G573, G621, G622, 
G776, G780, G784, G788, G812, G832, G836, G1509, G1517, G1525, 
G1533, G1581, G1621, G1629, G792, G796, G800, G804, G808, G816, 
G820, G824, G828, G871, G873, G875, G877, G879, G881, G883, 
G885, G1541, G1549, G1557, G1565, G1573, G1589, G1597, G1605, G1613, 
G1, G1513, G4, G1521, G7, G1529, G10, G1537, G28, G1585, 
G43, G1625, G46, G1633, G886, G2, G5, G8, G11, G13, 
G1545, G16, G1553, G19, G1561, G22, G1569, G25, G1577, G29, 
G31, G1593, G34, G1601, G37, G1609, G40, G1617, G44, G47, 
G857, G860, G863, G865, G14, G17, G20, G23, G26, G32, 
G35, G38, G41, G1913, G1921, G887, G462, G74, G1637, G1917, 
G1647, G1925, G1020, G1144, G1386, G1394, G1402, G1638, G1648, G1806, 
G1639, G1649, G287, G350, G427, G429, G431, G1028, G1152, G1392, 
G1400, G1408, G1812, G1216, G286, G349, G426, G428, G430, G67, 
G1643, G70, G1653, G1215, G49, G53, G59, G61, G65, G68, 
G71, G1217, G375, G1221, G376, G55;

not g0(G149, G101);
not g1(G153, G104);
not g2(G156, G107);
not g3(G160, G110);
not g4(G165, G113);
not g5(G168, G116);
not g6(G171, G119);
not g7(G175, G122);
not g8(G179, G125);
not g9(G184, G128);
not g10(G188, G131);
not g11(G191, G134);
not g12(G194, G137);
not g13(G198, G140);
not g14(G202, G143);
not g15(G206, G146);
nand g16(G231, G224, G898);
nand g17(G233, G227, G900);
not g18(G241, G237);
not g19(G244, G237);
assign G245 = G234;
assign G248 = G234;
not g22(G517, G469);
not g23(G529, G472);
not g24(G541, G475);
not g25(G553, G478);
not g26(G859, G953);
not g27(G862, G953);
not g28(G907, G898);
not g29(G909, G900);
assign G911 = G902;
not g31(G918, G902);
assign G919 = G902;
not g33(G922, G902);
assign G926 = G952;
not g35(G930, G952);
not g36(G932, G952);
assign G934 = G953;
not g38(G938, G953);
assign G943 = G953;
assign G947 = G953;
not g41(G949, G953);
assign G1506 = G101;
assign G1514 = G104;
assign G1522 = G107;
assign G1530 = G110;
assign G1538 = G113;
assign G1546 = G116;
assign G1554 = G119;
assign G1562 = G122;
assign G1570 = G125;
assign G1578 = G128;
assign G1586 = G131;
assign G1594 = G134;
assign G1602 = G137;
assign G1610 = G140;
assign G1618 = G143;
assign G1626 = G146;
not g58(G1512, G1506);
not g59(G1520, G1514);
not g60(G1528, G1522);
not g61(G1536, G1530);
not g62(G1544, G1538);
not g63(G1552, G1546);
not g64(G1560, G1554);
not g65(G1568, G1562);
not g66(G1576, G1570);
not g67(G1584, G1578);
not g68(G1592, G1586);
not g69(G1600, G1594);
not g70(G1608, G1602);
not g71(G1616, G1610);
not g72(G1624, G1618);
not g73(G1632, G1626);
nand g74(G50, G930, G947);
nand g75(G52, G930, G947);
nand g76(G56, G930, G947);
nand g77(G58, G930, G947);
nand g78(G62, G930, G947);
nand g79(G64, G930, G947);
assign G251 = G149;
assign G254 = G153;
assign G288 = G165;
assign G291 = G168;
assign G299 = G184;
assign G302 = G202;
and g86(G318, G224, G938);
assign G321 = G179;
assign G327 = G188;
assign G330 = G191;
and g90(G352, G227, G938);
assign G355 = G198;
and g92(G369, G210, G241, G938);
assign G382 = G206;
assign G385 = G198;
nand g95(G853, G943, G907);
nand g96(G856, G943, G909);
nand g97(G893, G248, G237);
nand g98(G954, G248, G922);
nand g99(G955, G244, G922);
assign G1050 = G160;
assign G1053 = G175;
assign G1176 = G179;
assign G1179 = G198;
assign G1197 = G149;
assign G1207 = G149;
assign G1222 = G153;
assign G1244 = G188;
assign G1278 = G156;
and g109(G1290, G217, G245, G938);
assign G1300 = G191;
assign G1312 = G160;
assign G1332 = G194;
and g113(G1335, G221, G245, G938);
assign G1442 = G517;
assign G1450 = G517;
assign G1458 = G529;
assign G1466 = G529;
assign G1474 = G541;
assign G1482 = G541;
assign G1490 = G553;
assign G1498 = G553;
and g122(G1634, G231, G934);
and g123(G1644, G233, G934);
assign G1657 = G156;
assign G1665 = G156;
assign G1697 = G171;
assign G1705 = G171;
assign G1713 = G206;
assign G1721 = G206;
assign G1745 = G194;
assign G1753 = G194;
assign G1785 = G160;
assign G1793 = G160;
assign G1814 = G165;
assign G1817 = G175;
and g136(G1830, G214, G241, G938);
assign G1833 = G202;
assign G1841 = G179;
assign G1849 = G179;
assign G1854 = G168;
assign G1857 = G175;
assign G1870 = G184;
assign G1873 = G202;
assign G1878 = G171;
assign G1881 = G184;
not g146(G1642, G1634);
not g147(G1652, G1644);
not g148(G1056, G1050);
not g149(G1057, G1053);
not g150(G1182, G1176);
not g151(G1183, G1179);
not g152(G1211, G1207);
not g153(G1298, G1290);
not g154(G1320, G1312);
not g155(G1338, G1332);
not g156(G1339, G1335);
and g157(G457, G210, G955);
and g158(G459, G217, G954);
nand g159(G482, G214, G955);
nand g160(G487, G221, G954);
nand g161(G492, G210, G955);
nand g162(G505, G217, G954);
not g163(G1456, G1450);
not g164(G1448, G1442);
not g165(G1472, G1466);
not g166(G1464, G1458);
not g167(G1488, G1482);
not g168(G1480, G1474);
not g169(G1504, G1498);
not g170(G1496, G1490);
nand g171(G956, G907, G919, G943, G893);
nand g172(G967, G909, G919, G943, G893);
nand g173(G978, G926, G949, G893);
and g174(G979, G926, G949, G893);
assign G980 = G251;
not g176(G1661, G1657);
assign G990 = G251;
not g178(G1669, G1665);
assign G1030 = G288;
not g180(G1701, G1697);
assign G1040 = G288;
not g182(G1709, G1705);
assign G1058 = G299;
not g184(G1717, G1713);
assign G1068 = G299;
not g186(G1725, G1721);
assign G1078 = G318;
assign G1090 = G318;
assign G1100 = G327;
not g190(G1749, G1745);
assign G1112 = G327;
not g192(G1757, G1753);
assign G1154 = G352;
not g194(G1789, G1785);
assign G1166 = G352;
not g196(G1797, G1793);
assign G1194 = G369;
not g198(G1201, G1197);
assign G1204 = G369;
not g200(G1820, G1814);
not g201(G1821, G1817);
not g202(G1230, G1222);
not g203(G1836, G1830);
not g204(G1837, G1833);
not g205(G1252, G1244);
assign G1256 = G382;
not g207(G1845, G1841);
assign G1268 = G382;
not g209(G1853, G1849);
not g210(G1860, G1854);
not g211(G1861, G1857);
not g212(G1286, G1278);
not g213(G1876, G1870);
not g214(G1877, G1873);
not g215(G1308, G1300);
not g216(G1884, G1878);
not g217(G1885, G1881);
assign G1654 = G254;
assign G1662 = G254;
assign G1694 = G291;
assign G1702 = G291;
assign G1710 = G302;
assign G1718 = G302;
assign G1726 = G321;
assign G1734 = G321;
assign G1742 = G330;
assign G1750 = G330;
assign G1782 = G355;
assign G1790 = G355;
assign G1838 = G385;
assign G1846 = G385;
nand g232(G297, G1053, G1056);
nand g233(G298, G1050, G1057);
nand g234(G361, G1179, G1182);
nand g235(G362, G1176, G1183);
nand g236(G404, G1335, G1338);
nand g237(G405, G1332, G1339);
nand g238(G1225, G1817, G1820);
nand g239(G1226, G1814, G1821);
nand g240(G1247, G1833, G1836);
nand g241(G1248, G1830, G1837);
nand g242(G1281, G1857, G1860);
nand g243(G1282, G1854, G1861);
nand g244(G1303, G1873, G1876);
nand g245(G1304, G1870, G1877);
nand g246(G1315, G1881, G1884);
nand g247(G1316, G1878, G1885);
not g248(G998, G990);
not g249(G988, G980);
nand g250(G268, G297, G298);
not g251(G1038, G1030);
not g252(G1048, G1040);
not g253(G1076, G1068);
not g254(G1066, G1058);
not g255(G1098, G1090);
not g256(G1120, G1112);
not g257(G1174, G1166);
nand g258(G363, G361, G362);
not g259(G1210, G1204);
nand g260(G373, G1204, G1211);
not g261(G1276, G1268);
nand g262(G406, G404, G405);
not g263(G565, G482);
assign G566 = G482;
not g265(G614, G487);
assign G615 = G487;
nand g267(G958, G956, G978);
nand g268(G969, G967, G978);
not g269(G1660, G1654);
nand g270(G984, G1654, G1661);
not g271(G1668, G1662);
nand g272(G994, G1662, G1669);
not g273(G1700, G1694);
nand g274(G1034, G1694, G1701);
not g275(G1708, G1702);
nand g276(G1044, G1702, G1709);
not g277(G1716, G1710);
nand g278(G1062, G1710, G1717);
not g279(G1724, G1718);
nand g280(G1072, G1718, G1725);
not g281(G1732, G1726);
not g282(G1086, G1078);
not g283(G1740, G1734);
not g284(G1748, G1742);
nand g285(G1104, G1742, G1749);
not g286(G1108, G1100);
not g287(G1756, G1750);
nand g288(G1116, G1750, G1757);
not g289(G1788, G1782);
nand g290(G1158, G1782, G1789);
not g291(G1162, G1154);
not g292(G1796, G1790);
nand g293(G1170, G1790, G1797);
not g294(G1200, G1194);
nand g295(G1203, G1194, G1201);
nand g296(G1227, G1225, G1226);
nand g297(G1249, G1247, G1248);
not g298(G1844, G1838);
nand g299(G1260, G1838, G1845);
not g300(G1264, G1256);
not g301(G1852, G1846);
nand g302(G1272, G1846, G1853);
nand g303(G1283, G1281, G1282);
nand g304(G1305, G1303, G1304);
nand g305(G1317, G1315, G1316);
assign G1410 = G492;
assign G1418 = G492;
assign G1426 = G505;
assign G1434 = G505;
not g310(G269, G268);
nand g311(G372, G1207, G1210);
nand g312(G983, G1657, G1660);
nand g313(G993, G1665, G1668);
nand g314(G1033, G1697, G1700);
nand g315(G1043, G1705, G1708);
nand g316(G1061, G1713, G1716);
nand g317(G1071, G1721, G1724);
nand g318(G1103, G1745, G1748);
nand g319(G1115, G1753, G1756);
nand g320(G1157, G1785, G1788);
nand g321(G1169, G1793, G1796);
not g322(G1184, G363);
nand g323(G1202, G1197, G1200);
nand g324(G1259, G1841, G1844);
nand g325(G1271, G1849, G1852);
not g326(G1322, G406);
nand g327(G374, G372, G373);
nand g328(G396, G1317, G1320);
not g329(G1321, G1317);
not g330(G1424, G1418);
not g331(G1416, G1410);
not g332(G1440, G1434);
not g333(G1432, G1426);
nand g334(G985, G983, G984);
nand g335(G995, G993, G994);
nand g336(G1035, G1033, G1034);
nand g337(G1045, G1043, G1044);
nand g338(G1063, G1061, G1062);
nand g339(G1073, G1071, G1072);
nand g340(G1105, G1103, G1104);
nand g341(G1117, G1115, G1116);
nand g342(G1159, G1157, G1158);
nand g343(G1171, G1169, G1170);
nand g344(G1212, G1202, G1203);
not g345(G1231, G1227);
nand g346(G1232, G1227, G1230);
not g347(G1253, G1249);
nand g348(G1254, G1249, G1252);
nand g349(G1261, G1259, G1260);
nand g350(G1273, G1271, G1272);
not g351(G1287, G1283);
nand g352(G1288, G1283, G1286);
not g353(G1309, G1305);
nand g354(G1310, G1305, G1308);
not g355(G1192, G1184);
nand g356(G397, G1312, G1321);
not g357(G1330, G1322);
assign G1000 = G269;
assign G1010 = G269;
nand g360(G1233, G1222, G1231);
nand g361(G1255, G1244, G1253);
nand g362(G1289, G1278, G1287);
nand g363(G1311, G1300, G1309);
not g364(G1381, G374);
nand g365(G257, G995, G998);
not g366(G999, G995);
nand g367(G260, G985, G988);
not g368(G989, G985);
nand g369(G272, G1035, G1038);
not g370(G1039, G1035);
nand g371(G294, G1045, G1048);
not g372(G1049, G1045);
nand g373(G305, G1073, G1076);
not g374(G1077, G1073);
nand g375(G308, G1063, G1066);
not g376(G1067, G1063);
nand g377(G333, G1117, G1120);
not g378(G1121, G1117);
nand g379(G358, G1171, G1174);
not g380(G1175, G1171);
not g381(G1220, G1212);
nand g382(G388, G1273, G1276);
not g383(G1277, G1273);
nand g384(G398, G396, G397);
not g385(G1109, G1105);
nand g386(G1110, G1105, G1108);
not g387(G1163, G1159);
nand g388(G1164, G1159, G1162);
nand g389(G1234, G1232, G1233);
not g390(G1265, G1261);
nand g391(G1266, G1261, G1264);
nand g392(G1822, G1254, G1255);
nand g393(G1862, G1310, G1311);
nand g394(G1865, G1288, G1289);
nand g395(G258, G990, G999);
nand g396(G261, G980, G989);
nand g397(G273, G1030, G1039);
not g398(G1018, G1010);
not g399(G1008, G1000);
nand g400(G295, G1040, G1049);
nand g401(G306, G1068, G1077);
nand g402(G309, G1058, G1067);
nand g403(G334, G1112, G1121);
nand g404(G359, G1166, G1175);
nand g405(G389, G1268, G1277);
not g406(G1385, G1381);
nand g407(G1111, G1100, G1109);
nand g408(G1165, G1154, G1163);
nand g409(G1267, G1256, G1265);
not g410(G1886, G398);
nand g411(G259, G257, G258);
nand g412(G262, G260, G261);
nand g413(G274, G272, G273);
nand g414(G296, G294, G295);
nand g415(G307, G305, G306);
nand g416(G310, G308, G309);
nand g417(G335, G333, G334);
nand g418(G360, G358, G359);
not g419(G1242, G1234);
nand g420(G390, G388, G389);
not g421(G1828, G1822);
not g422(G1868, G1862);
not g423(G1869, G1865);
nand g424(G1373, G1164, G1165);
nand g425(G1798, G1110, G1111);
nand g426(G1825, G1266, G1267);
not g427(G265, G259);
not g428(G314, G307);
not g429(G336, G335);
not g430(G407, G296);
nand g431(G1293, G1865, G1868);
nand g432(G1294, G1862, G1869);
not g433(G1892, G1886);
not g434(G1777, G360);
not g435(G1889, G390);
assign G410 = G310;
not g437(G1377, G1373);
not g438(G1804, G1798);
nand g439(G1237, G1825, G1828);
not g440(G1829, G1825);
nand g441(G1295, G1293, G1294);
assign G1670 = G274;
assign G1678 = G274;
assign G1729 = G310;
assign G1737 = G310;
assign G1761 = G262;
assign G1769 = G262;
assign G340 = G336;
assign G343 = G314;
not g450(G1781, G1777);
nand g451(G1238, G1822, G1829);
nand g452(G1325, G1889, G1892);
not g453(G1893, G1889);
assign G1340 = G407;
assign G1352 = G407;
assign G1673 = G265;
assign G1681 = G265;
assign G1801 = G314;
assign G1897 = G336;
assign G1905 = G336;
nand g461(G391, G1295, G1298);
not g462(G1299, G1295);
not g463(G1676, G1670);
not g464(G1684, G1678);
nand g465(G1081, G1729, G1732);
not g466(G1733, G1729);
nand g467(G1093, G1737, G1740);
not g468(G1741, G1737);
not g469(G1765, G1761);
not g470(G1773, G1769);
nand g471(G1239, G1237, G1238);
nand g472(G1326, G1886, G1893);
assign G1894 = G410;
assign G1902 = G410;
nand g475(G392, G1290, G1299);
not g476(G1360, G1352);
nand g477(G1003, G1673, G1676);
not g478(G1677, G1673);
nand g479(G1013, G1681, G1684);
not g480(G1685, G1681);
nand g481(G1082, G1726, G1733);
nand g482(G1094, G1734, G1741);
assign G1122 = G340;
assign G1134 = G340;
nand g485(G1187, G1801, G1804);
not g486(G1805, G1801);
nand g487(G1327, G1325, G1326);
not g488(G1901, G1897);
not g489(G1348, G1340);
not g490(G1909, G1905);
assign G1758 = G343;
assign G1766 = G343;
nand g493(G377, G1239, G1242);
not g494(G1243, G1239);
nand g495(G393, G391, G392);
nand g496(G1004, G1670, G1677);
nand g497(G1014, G1678, G1685);
nand g498(G1083, G1081, G1082);
nand g499(G1095, G1093, G1094);
nand g500(G1188, G1798, G1805);
not g501(G1900, G1894);
nand g502(G1344, G1894, G1901);
not g503(G1908, G1902);
nand g504(G1356, G1902, G1909);
not g505(G1142, G1134);
nand g506(G378, G1234, G1243);
nand g507(G399, G1327, G1330);
not g508(G1331, G1327);
nand g509(G1005, G1003, G1004);
nand g510(G1015, G1013, G1014);
not g511(G1764, G1758);
nand g512(G1126, G1758, G1765);
not g513(G1130, G1122);
not g514(G1772, G1766);
nand g515(G1138, G1766, G1773);
nand g516(G1189, G1187, G1188);
nand g517(G1343, G1897, G1900);
nand g518(G1355, G1905, G1908);
nand g519(G324, G1095, G1098);
not g520(G1099, G1095);
nand g521(G379, G377, G378);
nand g522(G400, G1322, G1331);
nand g523(G449, G393, G918);
not g524(G1087, G1083);
nand g525(G1088, G1083, G1086);
nand g526(G1125, G1761, G1764);
nand g527(G1137, G1769, G1772);
nand g528(G1345, G1343, G1344);
nand g529(G1357, G1355, G1356);
assign G1397 = G393;
nand g531(G277, G1015, G1018);
not g532(G1019, G1015);
nand g533(G280, G1005, G1008);
not g534(G1009, G1005);
nand g535(G325, G1090, G1099);
nand g536(G364, G1189, G1192);
not g537(G1193, G1189);
nand g538(G401, G399, G400);
nand g539(G1089, G1078, G1087);
nand g540(G1127, G1125, G1126);
nand g541(G1139, G1137, G1138);
nand g542(G278, G1010, G1019);
nand g543(G281, G1000, G1009);
nand g544(G326, G324, G325);
nand g545(G365, G1184, G1193);
nand g546(G413, G1357, G1360);
not g547(G1361, G1357);
not g548(G1401, G1397);
nand g549(G445, G379, G918);
not g550(G1349, G1345);
nand g551(G1350, G1345, G1348);
assign G1389 = G379;
assign G1493 = G449;
assign G1501 = G449;
nand g555(G1689, G1088, G1089);
nand g556(G279, G277, G278);
nand g557(G282, G280, G281);
nand g558(G346, G1139, G1142);
not g559(G1143, G1139);
nand g560(G366, G364, G365);
nand g561(G414, G1352, G1361);
nand g562(G453, G401, G918);
not g563(G1131, G1127);
nand g564(G1132, G1127, G1130);
nand g565(G1351, G1340, G1349);
not g566(G1365, G326);
assign G1405 = G401;
not g568(G285, G279);
nand g569(G347, G1134, G1143);
not g570(G367, G366);
nand g571(G415, G413, G414);
not g572(G1393, G1389);
nand g573(G556, G1501, G1504);
not g574(G1505, G1501);
nand g575(G559, G1493, G1496);
not g576(G1497, G1493);
not g577(G1693, G1689);
nand g578(G1133, G1122, G1131);
assign G1477 = G445;
assign G1485 = G445;
nand g581(G1809, G1350, G1351);
nand g582(G348, G346, G347);
not g583(G1369, G1365);
not g584(G1409, G1405);
nand g585(G557, G1498, G1505);
nand g586(G560, G1490, G1497);
assign G1362 = G282;
not g588(G1378, G415);
assign G1429 = G453;
assign G1437 = G453;
assign G1686 = G282;
nand g592(G1774, G1132, G1133);
and g593(G1910, G285, G853);
and g594(G1918, G856, G367);
nand g595(G544, G1485, G1488);
not g596(G1489, G1485);
nand g597(G547, G1477, G1480);
not g598(G1481, G1477);
nand g599(G558, G556, G557);
nand g600(G561, G559, G560);
not g601(G1813, G1809);
not g602(G1370, G348);
not g603(G1368, G1362);
nand g604(G417, G1362, G1369);
not g605(G1384, G1378);
nand g606(G424, G1378, G1385);
nand g607(G508, G1437, G1440);
not g608(G1441, G1437);
nand g609(G511, G1429, G1432);
not g610(G1433, G1429);
nand g611(G545, G1482, G1489);
nand g612(G548, G1474, G1481);
not g613(G564, G558);
not g614(G1692, G1686);
nand g615(G1024, G1686, G1693);
not g616(G1780, G1774);
nand g617(G1148, G1774, G1781);
not g618(G1916, G1910);
not g619(G1924, G1918);
nand g620(G416, G1365, G1368);
not g621(G1376, G1370);
nand g622(G421, G1370, G1377);
nand g623(G423, G1381, G1384);
nand g624(G509, G1434, G1441);
nand g625(G512, G1426, G1433);
nand g626(G546, G544, G545);
nand g627(G549, G547, G548);
not g628(G719, G561);
assign G722 = G561;
nand g630(G1023, G1689, G1692);
nand g631(G1147, G1777, G1780);
nand g632(G418, G416, G417);
nand g633(G420, G1373, G1376);
nand g634(G425, G423, G424);
nand g635(G510, G508, G509);
nand g636(G513, G511, G512);
not g637(G552, G546);
nand g638(G1025, G1023, G1024);
nand g639(G1149, G1147, G1148);
not g640(G419, G418);
nand g641(G422, G420, G421);
nand g642(G441, G425, G918);
not g643(G516, G510);
not g644(G725, G549);
assign G728 = G549;
not g646(G1029, G1025);
not g647(G1153, G1149);
nand g648(G433, G419, G918);
nand g649(G437, G422, G918);
not g650(G663, G513);
assign G666 = G513;
and g652(G731, G719, G725);
and g653(G746, G722, G725);
and g654(G756, G719, G728);
and g655(G770, G722, G728);
assign G1461 = G441;
assign G1469 = G441;
assign G1413 = G433;
assign G1421 = G433;
assign G1445 = G437;
assign G1453 = G437;
nand g662(G532, G1469, G1472);
not g663(G1473, G1469);
nand g664(G535, G1461, G1464);
not g665(G1465, G1461);
nand g666(G495, G1421, G1424);
not g667(G1425, G1421);
nand g668(G498, G1413, G1416);
not g669(G1417, G1413);
nand g670(G520, G1453, G1456);
not g671(G1457, G1453);
nand g672(G523, G1445, G1448);
not g673(G1449, G1445);
nand g674(G533, G1466, G1473);
nand g675(G536, G1458, G1465);
nand g676(G496, G1418, G1425);
nand g677(G499, G1410, G1417);
nand g678(G521, G1450, G1457);
nand g679(G524, G1442, G1449);
nand g680(G534, G532, G533);
nand g681(G537, G535, G536);
nand g682(G497, G495, G496);
nand g683(G500, G498, G499);
nand g684(G522, G520, G521);
nand g685(G525, G523, G524);
not g686(G540, G534);
not g687(G503, G497);
not g688(G528, G522);
not g689(G669, G537);
assign G672 = G537;
not g691(G569, G500);
and g692(G588, G566, G500);
not g693(G618, G525);
and g694(G639, G615, G525);
nand g695(G867, G516, G564, G552, G540, G482, G528, G503, G487);
assign G588a = G588;
assign G588b = G588;
assign G639a = G639;
assign G639b = G639;
and g700(G675, G663, G669);
and g701(G688, G666, G669);
and g702(G696, G663, G672);
and g703(G710, G666, G672);
and g704(G73, G949, G867, G932, G932);
and g705(G572, G565, G569);
and g706(G573, G566, G569);
and g707(G621, G614, G618);
and g708(G622, G615, G618);
nand g709(G776, G588a, G639a, G696, G731, G958);
nand g710(G780, G588a, G639a, G675, G756, G958);
nand g711(G784, G588a, G639a, G675, G746, G958);
nand g712(G788, G588a, G639a, G688, G731, G958);
nand g713(G812, G588b, G639a, G710, G746, G969);
nand g714(G832, G588b, G639b, G696, G770, G969);
nand g715(G836, G588b, G639b, G710, G756, G969);
and g716(G1509, G588a, G639a, G696, G731, G958);
and g717(G1517, G588a, G639a, G675, G756, G958);
and g718(G1525, G588a, G639a, G675, G746, G958);
and g719(G1533, G588a, G639a, G688, G731, G958);
and g720(G1581, G588b, G639a, G710, G746, G969);
and g721(G1621, G588b, G639b, G696, G770, G969);
and g722(G1629, G588b, G639b, G710, G756, G969);
nand g723(G792, G588a, G622, G696, G756, G958);
nand g724(G796, G588b, G622, G696, G746, G958);
nand g725(G800, G588b, G622, G710, G731, G958);
nand g726(G804, G588b, G622, G675, G770, G958);
nand g727(G808, G588b, G622, G688, G756, G969);
nand g728(G816, G573, G639b, G696, G756, G969);
nand g729(G820, G573, G639b, G696, G746, G969);
nand g730(G824, G573, G639b, G710, G731, G969);
nand g731(G828, G573, G639b, G688, G756, G969);
nand g732(G871, G588b, G622, G675, G731, G979);
nand g733(G873, G573, G639b, G675, G731, G979);
nand g734(G875, G573, G622, G696, G731, G979);
nand g735(G877, G573, G622, G675, G756, G979);
nand g736(G879, G573, G622, G675, G746, G979);
nand g737(G881, G573, G622, G688, G731, G979);
nand g738(G883, G573, G621, G675, G731, G979);
nand g739(G885, G572, G622, G675, G731, G979);
and g740(G1541, G588a, G622, G696, G756, G958);
and g741(G1549, G588b, G622, G696, G746, G958);
and g742(G1557, G588b, G622, G710, G731, G958);
and g743(G1565, G588b, G622, G675, G770, G958);
and g744(G1573, G588b, G622, G688, G756, G969);
and g745(G1589, G573, G639b, G696, G756, G969);
and g746(G1597, G573, G639b, G696, G746, G969);
and g747(G1605, G573, G639b, G710, G731, G969);
and g748(G1613, G573, G639b, G688, G756, G969);
nand g749(G1, G1509, G1512);
not g750(G1513, G1509);
nand g751(G4, G1517, G1520);
not g752(G1521, G1517);
nand g753(G7, G1525, G1528);
not g754(G1529, G1525);
nand g755(G10, G1533, G1536);
not g756(G1537, G1533);
nand g757(G28, G1581, G1584);
not g758(G1585, G1581);
nand g759(G43, G1621, G1624);
not g760(G1625, G1621);
nand g761(G46, G1629, G1632);
not g762(G1633, G1629);
and g763(G886, G871, G873, G875, G877, G879, G881, G883, G885);
nand g764(G2, G1506, G1513);
nand g765(G5, G1514, G1521);
nand g766(G8, G1522, G1529);
nand g767(G11, G1530, G1537);
nand g768(G13, G1541, G1544);
not g769(G1545, G1541);
nand g770(G16, G1549, G1552);
not g771(G1553, G1549);
nand g772(G19, G1557, G1560);
not g773(G1561, G1557);
nand g774(G22, G1565, G1568);
not g775(G1569, G1565);
nand g776(G25, G1573, G1576);
not g777(G1577, G1573);
nand g778(G29, G1578, G1585);
nand g779(G31, G1589, G1592);
not g780(G1593, G1589);
nand g781(G34, G1597, G1600);
not g782(G1601, G1597);
nand g783(G37, G1605, G1608);
not g784(G1609, G1605);
nand g785(G40, G1613, G1616);
not g786(G1617, G1613);
nand g787(G44, G1618, G1625);
nand g788(G47, G1626, G1633);
nand g789(G857, G776, G780, G784, G788, G792, G796, G800, G804);
nand g790(G860, G808, G812, G816, G820, G824, G828, G832, G836);
and g791(G863, G776, G780, G784, G788, G792, G796, G800, G804);
and g792(G865, G808, G812, G816, G820, G824, G828, G832, G836);
nand g793(G3, G1, G2);
nand g794(G6, G4, G5);
nand g795(G9, G7, G8);
nand g796(G12, G10, G11);
nand g797(G14, G1538, G1545);
nand g798(G17, G1546, G1553);
nand g799(G20, G1554, G1561);
nand g800(G23, G1562, G1569);
nand g801(G26, G1570, G1577);
nand g802(G30, G28, G29);
nand g803(G32, G1586, G1593);
nand g804(G35, G1594, G1601);
nand g805(G38, G1602, G1609);
nand g806(G41, G1610, G1617);
nand g807(G45, G43, G44);
nand g808(G48, G46, G47);
and g809(G1913, G857, G859);
and g810(G1921, G860, G862);
nand g811(G15, G13, G14);
nand g812(G18, G16, G17);
nand g813(G21, G19, G20);
nand g814(G24, G22, G23);
nand g815(G27, G25, G26);
nand g816(G33, G31, G32);
nand g817(G36, G34, G35);
nand g818(G39, G37, G38);
nand g819(G42, G40, G41);
and g820(G887, G863, G865, G886);
nand g821(G462, G863, G865);
and g822(G74, G949, G867, G952, G887);
nand g823(G1637, G1913, G1916);
not g824(G1917, G1913);
nand g825(G1647, G1921, G1924);
not g826(G1925, G1921);
nor g827(G75, G73, G74);
and g828(G1020, G457, G911, G462);
and g829(G1144, G469, G911, G462);
and g830(G1386, G475, G911, G462);
and g831(G1394, G478, G911, G462);
and g832(G1402, G459, G911, G462);
nand g833(G1638, G1910, G1917);
nand g834(G1648, G1918, G1925);
and g835(G1806, G472, G911, G462);
nand g836(G1639, G1637, G1638);
nand g837(G1649, G1647, G1648);
nand g838(G287, G1020, G1029);
nand g839(G350, G1144, G1153);
nand g840(G427, G1386, G1393);
nand g841(G429, G1394, G1401);
nand g842(G431, G1402, G1409);
not g843(G1028, G1020);
not g844(G1152, G1144);
not g845(G1392, G1386);
not g846(G1400, G1394);
not g847(G1408, G1402);
not g848(G1812, G1806);
nand g849(G1216, G1806, G1813);
nand g850(G286, G1025, G1028);
nand g851(G349, G1149, G1152);
nand g852(G426, G1389, G1392);
nand g853(G428, G1397, G1400);
nand g854(G430, G1405, G1408);
nand g855(G67, G1639, G1642);
not g856(G1643, G1639);
nand g857(G70, G1649, G1652);
not g858(G1653, G1649);
nand g859(G1215, G1809, G1812);
nand g860(G49, G286, G287);
nand g861(G53, G349, G350);
nand g862(G59, G426, G427);
nand g863(G61, G428, G429);
nand g864(G65, G430, G431);
nand g865(G68, G1634, G1643);
nand g866(G71, G1644, G1653);
nand g867(G1217, G1215, G1216);
and g868(G51, G49, G50);
and g869(G54, G52, G53);
and g870(G60, G58, G59);
and g871(G63, G61, G62);
and g872(G66, G64, G65);
nand g873(G69, G67, G68);
nand g874(G72, G70, G71);
nand g875(G375, G1217, G1220);
not g876(G1221, G1217);
nand g877(G376, G1212, G1221);
nand g878(G55, G375, G376);
and g879(G57, G55, G56);
endmodule
