
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729;

  XOR2X1 U429 ( .IN1(n397), .IN2(G32), .Q(G1355) );
  NAND2X0 U430 ( .IN1(n398), .IN2(n399), .QN(n397) );
  XOR2X1 U431 ( .IN1(n400), .IN2(G31), .Q(G1354) );
  NAND2X0 U432 ( .IN1(n398), .IN2(n401), .QN(n400) );
  XOR2X1 U433 ( .IN1(n402), .IN2(G30), .Q(G1353) );
  NAND2X0 U434 ( .IN1(n398), .IN2(n403), .QN(n402) );
  XOR2X1 U435 ( .IN1(n404), .IN2(G29), .Q(G1352) );
  NAND2X0 U436 ( .IN1(n398), .IN2(n405), .QN(n404) );
  AND4X1 U437 ( .IN1(n406), .IN2(n407), .IN3(n408), .IN4(n409), .Q(n398) );
  XNOR2X1 U438 ( .IN1(G28), .IN2(n410), .Q(G1351) );
  NOR2X0 U439 ( .IN1(n411), .IN2(n412), .QN(n410) );
  XNOR2X1 U440 ( .IN1(G27), .IN2(n413), .Q(G1350) );
  NOR2X0 U441 ( .IN1(n414), .IN2(n412), .QN(n413) );
  XNOR2X1 U442 ( .IN1(G26), .IN2(n415), .Q(G1349) );
  NOR2X0 U443 ( .IN1(n416), .IN2(n412), .QN(n415) );
  XNOR2X1 U444 ( .IN1(G25), .IN2(n417), .Q(G1348) );
  NOR2X0 U445 ( .IN1(n418), .IN2(n412), .QN(n417) );
  NAND4X0 U446 ( .IN1(n419), .IN2(n409), .IN3(n408), .IN4(n420), .QN(n412) );
  NOR2X0 U447 ( .IN1(n407), .IN2(n421), .QN(n420) );
  XNOR2X1 U448 ( .IN1(G24), .IN2(n422), .Q(G1347) );
  NOR2X0 U449 ( .IN1(n411), .IN2(n423), .QN(n422) );
  XNOR2X1 U450 ( .IN1(G23), .IN2(n424), .Q(G1346) );
  NOR2X0 U451 ( .IN1(n414), .IN2(n423), .QN(n424) );
  XNOR2X1 U452 ( .IN1(G22), .IN2(n425), .Q(G1345) );
  NOR2X0 U453 ( .IN1(n416), .IN2(n423), .QN(n425) );
  XNOR2X1 U454 ( .IN1(G21), .IN2(n426), .Q(G1344) );
  NOR2X0 U455 ( .IN1(n418), .IN2(n423), .QN(n426) );
  NAND4X0 U456 ( .IN1(n421), .IN2(n409), .IN3(n407), .IN4(n427), .QN(n423) );
  NOR2X0 U457 ( .IN1(n408), .IN2(n419), .QN(n427) );
  XOR2X1 U458 ( .IN1(n428), .IN2(G20), .Q(G1343) );
  NAND2X0 U459 ( .IN1(n429), .IN2(n399), .QN(n428) );
  XOR2X1 U460 ( .IN1(n430), .IN2(G19), .Q(G1342) );
  NAND2X0 U461 ( .IN1(n429), .IN2(n401), .QN(n430) );
  XNOR2X1 U462 ( .IN1(n431), .IN2(n432), .Q(G1341) );
  NAND2X0 U463 ( .IN1(n429), .IN2(n403), .QN(n431) );
  XOR2X1 U464 ( .IN1(n433), .IN2(G17), .Q(G1340) );
  NAND2X0 U465 ( .IN1(n429), .IN2(n405), .QN(n433) );
  AND4X1 U466 ( .IN1(n434), .IN2(n419), .IN3(n421), .IN4(n409), .Q(n429) );
  NAND2X0 U467 ( .IN1(n435), .IN2(n436), .QN(n409) );
  OR3X1 U468 ( .IN1(n403), .IN2(n437), .IN3(n399), .Q(n436) );
  OR3X1 U469 ( .IN1(n401), .IN2(n438), .IN3(n405), .Q(n435) );
  XOR2X1 U470 ( .IN1(n439), .IN2(G16), .Q(G1339) );
  NAND2X0 U471 ( .IN1(n440), .IN2(n441), .QN(n439) );
  XOR2X1 U472 ( .IN1(n442), .IN2(G15), .Q(G1338) );
  NAND2X0 U473 ( .IN1(n440), .IN2(n443), .QN(n442) );
  XOR2X1 U474 ( .IN1(n444), .IN2(G14), .Q(G1337) );
  NAND2X0 U475 ( .IN1(n440), .IN2(n445), .QN(n444) );
  XOR2X1 U476 ( .IN1(n446), .IN2(G13), .Q(G1336) );
  NAND2X0 U477 ( .IN1(n440), .IN2(n447), .QN(n446) );
  AND4X1 U478 ( .IN1(n438), .IN2(n418), .IN3(n414), .IN4(n448), .Q(n440) );
  NOR2X0 U479 ( .IN1(n416), .IN2(n411), .QN(n438) );
  XNOR2X1 U480 ( .IN1(G12), .IN2(n449), .Q(G1335) );
  NOR2X0 U481 ( .IN1(n419), .IN2(n450), .QN(n449) );
  XNOR2X1 U482 ( .IN1(G11), .IN2(n451), .Q(G1334) );
  NOR2X0 U483 ( .IN1(n407), .IN2(n450), .QN(n451) );
  XNOR2X1 U484 ( .IN1(G10), .IN2(n452), .Q(G1333) );
  NOR2X0 U485 ( .IN1(n421), .IN2(n450), .QN(n452) );
  XNOR2X1 U486 ( .IN1(G9), .IN2(n453), .Q(G1332) );
  NOR2X0 U487 ( .IN1(n408), .IN2(n450), .QN(n453) );
  NAND4X0 U488 ( .IN1(n418), .IN2(n448), .IN3(n411), .IN4(n454), .QN(n450) );
  NOR2X0 U489 ( .IN1(n414), .IN2(n416), .QN(n454) );
  XNOR2X1 U490 ( .IN1(G8), .IN2(n455), .Q(G1331) );
  NOR2X0 U491 ( .IN1(n419), .IN2(n456), .QN(n455) );
  XNOR2X1 U492 ( .IN1(G7), .IN2(n457), .Q(G1330) );
  NOR2X0 U493 ( .IN1(n407), .IN2(n456), .QN(n457) );
  XNOR2X1 U494 ( .IN1(G6), .IN2(n458), .Q(G1329) );
  NOR2X0 U495 ( .IN1(n421), .IN2(n456), .QN(n458) );
  XNOR2X1 U496 ( .IN1(G5), .IN2(n459), .Q(G1328) );
  NOR2X0 U497 ( .IN1(n408), .IN2(n456), .QN(n459) );
  NAND4X0 U498 ( .IN1(n414), .IN2(n448), .IN3(n416), .IN4(n460), .QN(n456) );
  NOR2X0 U499 ( .IN1(n411), .IN2(n418), .QN(n460) );
  XOR2X1 U500 ( .IN1(n461), .IN2(G4), .Q(G1327) );
  NAND2X0 U501 ( .IN1(n462), .IN2(n441), .QN(n461) );
  XOR2X1 U502 ( .IN1(n463), .IN2(G3), .Q(G1326) );
  NAND2X0 U503 ( .IN1(n462), .IN2(n443), .QN(n463) );
  XOR2X1 U504 ( .IN1(n464), .IN2(G2), .Q(G1325) );
  NAND2X0 U505 ( .IN1(n462), .IN2(n445), .QN(n464) );
  XOR2X1 U506 ( .IN1(n465), .IN2(G1), .Q(G1324) );
  NAND2X0 U507 ( .IN1(n462), .IN2(n447), .QN(n465) );
  AND4X1 U508 ( .IN1(n437), .IN2(n411), .IN3(n416), .IN4(n448), .Q(n462) );
  NAND2X0 U509 ( .IN1(n466), .IN2(n467), .QN(n448) );
  OR3X1 U510 ( .IN1(n445), .IN2(n434), .IN3(n441), .Q(n467) );
  NOR2X0 U511 ( .IN1(n408), .IN2(n407), .QN(n434) );
  INVX0 U512 ( .INP(n443), .ZN(n407) );
  INVX0 U513 ( .INP(n447), .ZN(n408) );
  OR3X1 U514 ( .IN1(n447), .IN2(n406), .IN3(n443), .Q(n466) );
  MUX21X1 U515 ( .IN1(n468), .IN2(n469), .S(n470), .Q(n443) );
  NOR2X0 U516 ( .IN1(n471), .IN2(n472), .QN(n470) );
  XOR2X1 U517 ( .IN1(keyinput68), .IN2(n473), .Q(n472) );
  AND2X1 U518 ( .IN1(n474), .IN2(n475), .Q(n473) );
  XOR2X1 U519 ( .IN1(n476), .IN2(keyinput69), .Q(n471) );
  NAND2X0 U520 ( .IN1(n475), .IN2(n477), .QN(n476) );
  XOR2X1 U521 ( .IN1(n478), .IN2(keyinput42), .Q(n475) );
  NAND2X0 U522 ( .IN1(n474), .IN2(n477), .QN(n478) );
  XNOR3X1 U523 ( .IN1(keyinput21), .IN2(G15), .IN3(G11), .Q(n477) );
  XNOR3X1 U524 ( .IN1(keyinput20), .IN2(G7), .IN3(G3), .Q(n474) );
  NOR2X0 U525 ( .IN1(n479), .IN2(n480), .QN(n469) );
  OR2X1 U526 ( .IN1(n480), .IN2(n479), .Q(n468) );
  AOI21X1 U527 ( .IN1(G35), .IN2(G41), .IN3(n481), .QN(n479) );
  XNOR2X1 U528 ( .IN1(n482), .IN2(keyinput122), .Q(n480) );
  NAND3X0 U529 ( .IN1(G41), .IN2(n481), .IN3(G35), .QN(n482) );
  XOR2X1 U530 ( .IN1(keyinput118), .IN2(n483), .Q(n481) );
  AND2X1 U531 ( .IN1(n484), .IN2(n485), .Q(n483) );
  XOR2X1 U532 ( .IN1(keyinput109), .IN2(n486), .Q(n485) );
  AND2X1 U533 ( .IN1(n487), .IN2(n488), .Q(n486) );
  XOR2X1 U534 ( .IN1(n489), .IN2(keyinput108), .Q(n484) );
  NAND2X0 U535 ( .IN1(n488), .IN2(n490), .QN(n489) );
  XOR2X1 U536 ( .IN1(n491), .IN2(keyinput94), .Q(n488) );
  NAND2X0 U537 ( .IN1(n490), .IN2(n487), .QN(n491) );
  NOR2X0 U538 ( .IN1(n421), .IN2(n419), .QN(n406) );
  INVX0 U539 ( .INP(n441), .ZN(n419) );
  MUX21X1 U540 ( .IN1(n492), .IN2(n493), .S(n494), .Q(n441) );
  NOR2X0 U541 ( .IN1(n495), .IN2(n496), .QN(n494) );
  XOR2X1 U542 ( .IN1(keyinput71), .IN2(n497), .Q(n496) );
  AND2X1 U543 ( .IN1(n498), .IN2(n499), .Q(n497) );
  XOR2X1 U544 ( .IN1(n500), .IN2(keyinput70), .Q(n495) );
  NAND2X0 U545 ( .IN1(n501), .IN2(n499), .QN(n500) );
  XNOR2X1 U546 ( .IN1(n502), .IN2(keyinput43), .Q(n499) );
  NAND2X0 U547 ( .IN1(n501), .IN2(n498), .QN(n502) );
  XOR3X1 U548 ( .IN1(keyinput23), .IN2(G16), .IN3(G12), .Q(n498) );
  XNOR3X1 U549 ( .IN1(keyinput22), .IN2(G8), .IN3(G4), .Q(n501) );
  NOR2X0 U550 ( .IN1(n503), .IN2(n504), .QN(n493) );
  OR2X1 U551 ( .IN1(n504), .IN2(n503), .Q(n492) );
  AOI21X1 U552 ( .IN1(G36), .IN2(G41), .IN3(n505), .QN(n503) );
  XNOR2X1 U553 ( .IN1(n506), .IN2(keyinput123), .Q(n504) );
  NAND3X0 U554 ( .IN1(G36), .IN2(G41), .IN3(n505), .QN(n506) );
  XOR2X1 U555 ( .IN1(n507), .IN2(keyinput119), .Q(n505) );
  NAND2X0 U556 ( .IN1(n508), .IN2(n509), .QN(n507) );
  XOR2X1 U557 ( .IN1(keyinput110), .IN2(n510), .Q(n509) );
  AND2X1 U558 ( .IN1(n511), .IN2(n512), .Q(n510) );
  XOR2X1 U559 ( .IN1(n513), .IN2(keyinput111), .Q(n508) );
  NAND2X0 U560 ( .IN1(n512), .IN2(n514), .QN(n513) );
  XOR2X1 U561 ( .IN1(n515), .IN2(keyinput95), .Q(n512) );
  NAND2X0 U562 ( .IN1(n511), .IN2(n514), .QN(n515) );
  INVX0 U563 ( .INP(n445), .ZN(n421) );
  MUX21X1 U564 ( .IN1(n516), .IN2(n517), .S(n518), .Q(n445) );
  NOR2X0 U565 ( .IN1(n519), .IN2(n520), .QN(n518) );
  XOR2X1 U566 ( .IN1(keyinput67), .IN2(n521), .Q(n520) );
  AND2X1 U567 ( .IN1(n522), .IN2(n523), .Q(n521) );
  XOR2X1 U568 ( .IN1(n524), .IN2(keyinput66), .Q(n519) );
  NAND2X0 U569 ( .IN1(n523), .IN2(n525), .QN(n524) );
  XNOR2X1 U570 ( .IN1(n526), .IN2(keyinput41), .Q(n523) );
  NAND2X0 U571 ( .IN1(n522), .IN2(n525), .QN(n526) );
  XOR3X1 U572 ( .IN1(keyinput18), .IN2(G6), .IN3(G2), .Q(n525) );
  XOR3X1 U573 ( .IN1(keyinput19), .IN2(G14), .IN3(G10), .Q(n522) );
  AND2X1 U574 ( .IN1(n527), .IN2(n528), .Q(n517) );
  NAND2X0 U575 ( .IN1(n528), .IN2(n527), .QN(n516) );
  AO21X1 U576 ( .IN1(G34), .IN2(G41), .IN3(n529), .Q(n527) );
  XNOR2X1 U577 ( .IN1(n530), .IN2(keyinput121), .Q(n528) );
  NAND3X0 U578 ( .IN1(G34), .IN2(G41), .IN3(n529), .QN(n530) );
  XOR2X1 U579 ( .IN1(n531), .IN2(keyinput117), .Q(n529) );
  NAND2X0 U580 ( .IN1(n532), .IN2(n533), .QN(n531) );
  XOR2X1 U581 ( .IN1(keyinput106), .IN2(n534), .Q(n533) );
  AND2X1 U582 ( .IN1(n487), .IN2(n535), .Q(n534) );
  XOR2X1 U583 ( .IN1(n536), .IN2(keyinput107), .Q(n532) );
  NAND2X0 U584 ( .IN1(n535), .IN2(n514), .QN(n536) );
  XOR2X1 U585 ( .IN1(n537), .IN2(keyinput93), .Q(n535) );
  NAND2X0 U586 ( .IN1(n487), .IN2(n514), .QN(n537) );
  XNOR2X1 U587 ( .IN1(n538), .IN2(keyinput87), .Q(n514) );
  NAND2X0 U588 ( .IN1(n539), .IN2(n540), .QN(n538) );
  XOR2X1 U589 ( .IN1(keyinput63), .IN2(n541), .Q(n540) );
  AND2X1 U590 ( .IN1(n542), .IN2(n543), .Q(n541) );
  XOR2X1 U591 ( .IN1(n544), .IN2(keyinput62), .Q(n539) );
  NAND2X0 U592 ( .IN1(n545), .IN2(n543), .QN(n544) );
  XNOR2X1 U593 ( .IN1(n546), .IN2(keyinput39), .Q(n543) );
  NAND2X0 U594 ( .IN1(n545), .IN2(n542), .QN(n546) );
  XOR3X1 U595 ( .IN1(keyinput15), .IN2(G32), .IN3(G31), .Q(n542) );
  XNOR3X1 U596 ( .IN1(keyinput14), .IN2(G30), .IN3(G29), .Q(n545) );
  XOR2X1 U597 ( .IN1(n547), .IN2(keyinput86), .Q(n487) );
  NAND2X0 U598 ( .IN1(n548), .IN2(n549), .QN(n547) );
  XOR2X1 U599 ( .IN1(keyinput61), .IN2(n550), .Q(n549) );
  AND2X1 U600 ( .IN1(n551), .IN2(n552), .Q(n550) );
  XOR2X1 U601 ( .IN1(n553), .IN2(keyinput60), .Q(n548) );
  NAND2X0 U602 ( .IN1(n554), .IN2(n551), .QN(n553) );
  XNOR2X1 U603 ( .IN1(n555), .IN2(keyinput38), .Q(n551) );
  NAND2X0 U604 ( .IN1(n552), .IN2(n554), .QN(n555) );
  XNOR3X1 U605 ( .IN1(keyinput13), .IN2(G28), .IN3(G27), .Q(n552) );
  XNOR3X1 U606 ( .IN1(keyinput12), .IN2(G26), .IN3(G25), .Q(n554) );
  MUX21X1 U607 ( .IN1(n556), .IN2(n557), .S(n558), .Q(n447) );
  NOR2X0 U608 ( .IN1(n559), .IN2(n560), .QN(n558) );
  XOR2X1 U609 ( .IN1(keyinput65), .IN2(n561), .Q(n560) );
  NOR2X0 U610 ( .IN1(n562), .IN2(n563), .QN(n561) );
  XOR2X1 U611 ( .IN1(keyinput64), .IN2(n564), .Q(n559) );
  NOR2X0 U612 ( .IN1(n565), .IN2(n563), .QN(n564) );
  XNOR2X1 U613 ( .IN1(n566), .IN2(keyinput40), .Q(n563) );
  OR2X1 U614 ( .IN1(n565), .IN2(n562), .Q(n566) );
  XNOR3X1 U615 ( .IN1(keyinput17), .IN2(G9), .IN3(G13), .Q(n562) );
  XOR3X1 U616 ( .IN1(keyinput16), .IN2(G5), .IN3(G1), .Q(n565) );
  AND2X1 U617 ( .IN1(n567), .IN2(n568), .Q(n557) );
  NAND2X0 U618 ( .IN1(n568), .IN2(n567), .QN(n556) );
  AO21X1 U619 ( .IN1(G33), .IN2(G41), .IN3(n569), .Q(n567) );
  XNOR2X1 U620 ( .IN1(n570), .IN2(keyinput120), .Q(n568) );
  NAND3X0 U621 ( .IN1(G41), .IN2(n569), .IN3(G33), .QN(n570) );
  XOR2X1 U622 ( .IN1(keyinput116), .IN2(n571), .Q(n569) );
  AND2X1 U623 ( .IN1(n572), .IN2(n573), .Q(n571) );
  XOR2X1 U624 ( .IN1(keyinput105), .IN2(n574), .Q(n573) );
  AND2X1 U625 ( .IN1(n511), .IN2(n575), .Q(n574) );
  XOR2X1 U626 ( .IN1(n576), .IN2(keyinput104), .Q(n572) );
  NAND2X0 U627 ( .IN1(n575), .IN2(n490), .QN(n576) );
  XOR2X1 U628 ( .IN1(n577), .IN2(keyinput92), .Q(n575) );
  NAND2X0 U629 ( .IN1(n490), .IN2(n511), .QN(n577) );
  XNOR2X1 U630 ( .IN1(n578), .IN2(keyinput85), .Q(n511) );
  NAND2X0 U631 ( .IN1(n579), .IN2(n580), .QN(n578) );
  XOR2X1 U632 ( .IN1(keyinput58), .IN2(n581), .Q(n580) );
  NOR2X0 U633 ( .IN1(n582), .IN2(n583), .QN(n581) );
  XOR2X1 U634 ( .IN1(keyinput59), .IN2(n584), .Q(n579) );
  NOR2X0 U635 ( .IN1(n582), .IN2(n585), .QN(n584) );
  XOR2X1 U636 ( .IN1(n586), .IN2(keyinput37), .Q(n582) );
  OR2X1 U637 ( .IN1(n583), .IN2(n585), .Q(n586) );
  XOR3X1 U638 ( .IN1(keyinput11), .IN2(G24), .IN3(G23), .Q(n585) );
  XOR3X1 U639 ( .IN1(keyinput10), .IN2(G22), .IN3(G21), .Q(n583) );
  XOR2X1 U640 ( .IN1(n587), .IN2(keyinput84), .Q(n490) );
  NAND2X0 U641 ( .IN1(n588), .IN2(n589), .QN(n587) );
  XOR2X1 U642 ( .IN1(keyinput56), .IN2(n590), .Q(n589) );
  NOR2X0 U643 ( .IN1(n591), .IN2(n592), .QN(n590) );
  XOR2X1 U644 ( .IN1(keyinput57), .IN2(n593), .Q(n588) );
  NOR2X0 U645 ( .IN1(n594), .IN2(n592), .QN(n593) );
  XNOR2X1 U646 ( .IN1(n595), .IN2(keyinput36), .Q(n592) );
  OR2X1 U647 ( .IN1(n591), .IN2(n594), .Q(n595) );
  XNOR3X1 U648 ( .IN1(keyinput8), .IN2(n432), .IN3(G17), .Q(n591) );
  INVX0 U649 ( .INP(G18), .ZN(n432) );
  XNOR3X1 U650 ( .IN1(keyinput9), .IN2(G20), .IN3(G19), .Q(n594) );
  INVX0 U651 ( .INP(n403), .ZN(n416) );
  MUX21X1 U652 ( .IN1(n596), .IN2(n597), .S(n598), .Q(n403) );
  NOR2X0 U653 ( .IN1(n599), .IN2(n600), .QN(n598) );
  XOR2X1 U654 ( .IN1(n601), .IN2(keyinput75), .Q(n600) );
  NAND2X0 U655 ( .IN1(n602), .IN2(n603), .QN(n601) );
  XOR2X1 U656 ( .IN1(n604), .IN2(keyinput74), .Q(n599) );
  NAND2X0 U657 ( .IN1(n602), .IN2(n605), .QN(n604) );
  XOR2X1 U658 ( .IN1(n606), .IN2(keyinput45), .Q(n602) );
  NAND2X0 U659 ( .IN1(n605), .IN2(n603), .QN(n606) );
  XNOR3X1 U660 ( .IN1(keyinput27), .IN2(G30), .IN3(G26), .Q(n603) );
  XNOR3X1 U661 ( .IN1(keyinput26), .IN2(G22), .IN3(G18), .Q(n605) );
  NOR2X0 U662 ( .IN1(n607), .IN2(n608), .QN(n597) );
  OR2X1 U663 ( .IN1(n608), .IN2(n607), .Q(n596) );
  AOI21X1 U664 ( .IN1(G38), .IN2(G41), .IN3(n609), .QN(n607) );
  XNOR2X1 U665 ( .IN1(n610), .IN2(keyinput125), .Q(n608) );
  NAND3X0 U666 ( .IN1(G41), .IN2(n609), .IN3(G38), .QN(n610) );
  XOR2X1 U667 ( .IN1(keyinput113), .IN2(n611), .Q(n609) );
  AND2X1 U668 ( .IN1(n612), .IN2(n613), .Q(n611) );
  XOR2X1 U669 ( .IN1(keyinput99), .IN2(n614), .Q(n613) );
  NOR2X0 U670 ( .IN1(n615), .IN2(n616), .QN(n614) );
  XOR2X1 U671 ( .IN1(n617), .IN2(keyinput98), .Q(n612) );
  OR2X1 U672 ( .IN1(n616), .IN2(n618), .Q(n617) );
  XNOR2X1 U673 ( .IN1(n619), .IN2(keyinput89), .Q(n616) );
  NAND2X0 U674 ( .IN1(n620), .IN2(n621), .QN(n619) );
  INVX0 U675 ( .INP(n399), .ZN(n411) );
  MUX21X1 U676 ( .IN1(n622), .IN2(n623), .S(n624), .Q(n399) );
  NOR2X0 U677 ( .IN1(n625), .IN2(n626), .QN(n624) );
  XOR2X1 U678 ( .IN1(n627), .IN2(keyinput79), .Q(n626) );
  NAND2X0 U679 ( .IN1(n628), .IN2(n629), .QN(n627) );
  XOR2X1 U680 ( .IN1(n630), .IN2(keyinput78), .Q(n625) );
  NAND2X0 U681 ( .IN1(n628), .IN2(n631), .QN(n630) );
  XOR2X1 U682 ( .IN1(n632), .IN2(keyinput47), .Q(n628) );
  NAND2X0 U683 ( .IN1(n631), .IN2(n629), .QN(n632) );
  XNOR3X1 U684 ( .IN1(keyinput31), .IN2(G32), .IN3(G28), .Q(n629) );
  XNOR3X1 U685 ( .IN1(keyinput30), .IN2(G24), .IN3(G20), .Q(n631) );
  AND2X1 U686 ( .IN1(n633), .IN2(n634), .Q(n623) );
  NAND2X0 U687 ( .IN1(n634), .IN2(n633), .QN(n622) );
  AO21X1 U688 ( .IN1(G40), .IN2(G41), .IN3(n635), .Q(n633) );
  XNOR2X1 U689 ( .IN1(n636), .IN2(keyinput127), .Q(n634) );
  NAND3X0 U690 ( .IN1(G40), .IN2(G41), .IN3(n635), .QN(n636) );
  XOR2X1 U691 ( .IN1(n637), .IN2(keyinput115), .Q(n635) );
  NAND2X0 U692 ( .IN1(n638), .IN2(n639), .QN(n637) );
  XOR2X1 U693 ( .IN1(keyinput102), .IN2(n640), .Q(n639) );
  NOR2X0 U694 ( .IN1(n641), .IN2(n642), .QN(n640) );
  INVX0 U695 ( .INP(n643), .ZN(n641) );
  XOR2X1 U696 ( .IN1(keyinput103), .IN2(n644), .Q(n638) );
  NOR2X0 U697 ( .IN1(n642), .IN2(n615), .QN(n644) );
  XOR2X1 U698 ( .IN1(n645), .IN2(keyinput91), .Q(n642) );
  NAND2X0 U699 ( .IN1(n620), .IN2(n643), .QN(n645) );
  INVX0 U700 ( .INP(n615), .ZN(n620) );
  XNOR2X1 U701 ( .IN1(n646), .IN2(keyinput83), .Q(n615) );
  NAND2X0 U702 ( .IN1(n647), .IN2(n648), .QN(n646) );
  XOR2X1 U703 ( .IN1(keyinput55), .IN2(n649), .Q(n648) );
  AND2X1 U704 ( .IN1(n650), .IN2(n651), .Q(n649) );
  XOR2X1 U705 ( .IN1(n652), .IN2(keyinput54), .Q(n647) );
  NAND2X0 U706 ( .IN1(n653), .IN2(n651), .QN(n652) );
  XNOR2X1 U707 ( .IN1(n654), .IN2(keyinput35), .Q(n651) );
  NAND2X0 U708 ( .IN1(n653), .IN2(n650), .QN(n654) );
  XOR3X1 U709 ( .IN1(keyinput7), .IN2(G16), .IN3(G15), .Q(n650) );
  XNOR3X1 U710 ( .IN1(keyinput6), .IN2(G14), .IN3(G13), .Q(n653) );
  NOR2X0 U711 ( .IN1(n414), .IN2(n418), .QN(n437) );
  INVX0 U712 ( .INP(n405), .ZN(n418) );
  MUX21X1 U713 ( .IN1(n655), .IN2(n656), .S(n657), .Q(n405) );
  NOR2X0 U714 ( .IN1(n658), .IN2(n659), .QN(n657) );
  XOR2X1 U715 ( .IN1(keyinput73), .IN2(n660), .Q(n659) );
  AND2X1 U716 ( .IN1(n661), .IN2(n662), .Q(n660) );
  XOR2X1 U717 ( .IN1(n663), .IN2(keyinput72), .Q(n658) );
  NAND2X0 U718 ( .IN1(n662), .IN2(n664), .QN(n663) );
  XOR2X1 U719 ( .IN1(n665), .IN2(keyinput44), .Q(n662) );
  NAND2X0 U720 ( .IN1(n661), .IN2(n664), .QN(n665) );
  XOR3X1 U721 ( .IN1(keyinput24), .IN2(G21), .IN3(G17), .Q(n664) );
  XOR3X1 U722 ( .IN1(keyinput25), .IN2(G29), .IN3(G25), .Q(n661) );
  NOR2X0 U723 ( .IN1(n666), .IN2(n667), .QN(n656) );
  OR2X1 U724 ( .IN1(n667), .IN2(n666), .Q(n655) );
  AOI21X1 U725 ( .IN1(G37), .IN2(G41), .IN3(n668), .QN(n666) );
  XNOR2X1 U726 ( .IN1(n669), .IN2(keyinput124), .Q(n667) );
  NAND3X0 U727 ( .IN1(G37), .IN2(G41), .IN3(n668), .QN(n669) );
  XOR2X1 U728 ( .IN1(n670), .IN2(keyinput112), .Q(n668) );
  NAND2X0 U729 ( .IN1(n671), .IN2(n672), .QN(n670) );
  XOR2X1 U730 ( .IN1(keyinput96), .IN2(n673), .Q(n672) );
  AND2X1 U731 ( .IN1(n674), .IN2(n675), .Q(n673) );
  XOR2X1 U732 ( .IN1(n676), .IN2(keyinput97), .Q(n671) );
  NAND2X0 U733 ( .IN1(n674), .IN2(n643), .QN(n676) );
  XNOR2X1 U734 ( .IN1(n677), .IN2(keyinput88), .Q(n674) );
  NAND2X0 U735 ( .IN1(n675), .IN2(n643), .QN(n677) );
  XNOR2X1 U736 ( .IN1(n678), .IN2(keyinput81), .Q(n643) );
  NAND2X0 U737 ( .IN1(n679), .IN2(n680), .QN(n678) );
  XOR2X1 U738 ( .IN1(keyinput50), .IN2(n681), .Q(n680) );
  AND2X1 U739 ( .IN1(n682), .IN2(n683), .Q(n681) );
  XOR2X1 U740 ( .IN1(n684), .IN2(keyinput51), .Q(n679) );
  NAND2X0 U741 ( .IN1(n685), .IN2(n682), .QN(n684) );
  XNOR2X1 U742 ( .IN1(n686), .IN2(keyinput33), .Q(n682) );
  NAND2X0 U743 ( .IN1(n683), .IN2(n685), .QN(n686) );
  XNOR3X1 U744 ( .IN1(keyinput2), .IN2(G6), .IN3(G5), .Q(n683) );
  XNOR3X1 U745 ( .IN1(keyinput3), .IN2(G8), .IN3(G7), .Q(n685) );
  INVX0 U746 ( .INP(n401), .ZN(n414) );
  MUX21X1 U747 ( .IN1(n687), .IN2(n688), .S(n689), .Q(n401) );
  NOR2X0 U748 ( .IN1(n690), .IN2(n691), .QN(n689) );
  XOR2X1 U749 ( .IN1(keyinput76), .IN2(n692), .Q(n691) );
  AND2X1 U750 ( .IN1(n693), .IN2(n694), .Q(n692) );
  XOR2X1 U751 ( .IN1(n695), .IN2(keyinput77), .Q(n690) );
  NAND2X0 U752 ( .IN1(n694), .IN2(n696), .QN(n695) );
  XOR2X1 U753 ( .IN1(n697), .IN2(keyinput46), .Q(n694) );
  NAND2X0 U754 ( .IN1(n693), .IN2(n696), .QN(n697) );
  XOR3X1 U755 ( .IN1(keyinput29), .IN2(G31), .IN3(G27), .Q(n696) );
  XNOR3X1 U756 ( .IN1(keyinput28), .IN2(G23), .IN3(G19), .Q(n693) );
  AND2X1 U757 ( .IN1(n698), .IN2(n699), .Q(n688) );
  NAND2X0 U758 ( .IN1(n699), .IN2(n698), .QN(n687) );
  AO21X1 U759 ( .IN1(G41), .IN2(G39), .IN3(n700), .Q(n698) );
  XNOR2X1 U760 ( .IN1(n701), .IN2(keyinput126), .Q(n699) );
  NAND3X0 U761 ( .IN1(G39), .IN2(n700), .IN3(G41), .QN(n701) );
  XOR2X1 U762 ( .IN1(keyinput114), .IN2(n702), .Q(n700) );
  AND2X1 U763 ( .IN1(n703), .IN2(n704), .Q(n702) );
  XOR2X1 U764 ( .IN1(keyinput100), .IN2(n705), .Q(n704) );
  NOR2X0 U765 ( .IN1(n706), .IN2(n707), .QN(n705) );
  XOR2X1 U766 ( .IN1(keyinput101), .IN2(n708), .Q(n703) );
  NOR2X0 U767 ( .IN1(n618), .IN2(n707), .QN(n708) );
  XNOR2X1 U768 ( .IN1(n709), .IN2(keyinput90), .Q(n707) );
  NAND2X0 U769 ( .IN1(n675), .IN2(n621), .QN(n709) );
  INVX0 U770 ( .INP(n706), .ZN(n675) );
  XNOR2X1 U771 ( .IN1(n710), .IN2(keyinput80), .Q(n706) );
  NAND2X0 U772 ( .IN1(n711), .IN2(n712), .QN(n710) );
  XOR2X1 U773 ( .IN1(n713), .IN2(keyinput48), .Q(n712) );
  NAND2X0 U774 ( .IN1(n714), .IN2(n715), .QN(n713) );
  XOR2X1 U775 ( .IN1(n716), .IN2(keyinput49), .Q(n711) );
  NAND2X0 U776 ( .IN1(n714), .IN2(n717), .QN(n716) );
  XOR2X1 U777 ( .IN1(n718), .IN2(keyinput32), .Q(n714) );
  NAND2X0 U778 ( .IN1(n717), .IN2(n715), .QN(n718) );
  XOR3X1 U779 ( .IN1(keyinput0), .IN2(G2), .IN3(G1), .Q(n715) );
  XNOR3X1 U780 ( .IN1(keyinput1), .IN2(G4), .IN3(G3), .Q(n717) );
  INVX0 U781 ( .INP(n621), .ZN(n618) );
  XNOR2X1 U782 ( .IN1(n719), .IN2(keyinput82), .Q(n621) );
  NAND2X0 U783 ( .IN1(n720), .IN2(n721), .QN(n719) );
  XOR2X1 U784 ( .IN1(keyinput53), .IN2(n722), .Q(n721) );
  AND2X1 U785 ( .IN1(n723), .IN2(n724), .Q(n722) );
  XOR2X1 U786 ( .IN1(n725), .IN2(keyinput52), .Q(n720) );
  NAND2X0 U787 ( .IN1(n726), .IN2(n723), .QN(n725) );
  XNOR2X1 U788 ( .IN1(n727), .IN2(keyinput34), .Q(n723) );
  NAND2X0 U789 ( .IN1(n724), .IN2(n726), .QN(n727) );
  XNOR3X1 U790 ( .IN1(keyinput5), .IN2(G12), .IN3(G11), .Q(n724) );
  XNOR3X1 U791 ( .IN1(keyinput4), .IN2(n728), .IN3(n729), .Q(n726) );
  INVX0 U792 ( .INP(G10), .ZN(n729) );
  INVX0 U793 ( .INP(G9), .ZN(n728) );
endmodule

