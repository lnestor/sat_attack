
module c499 ( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, 
        N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, 
        N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, 
        N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, 
        N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, 
        N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, keyinput0, 
        keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, 
        keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, 
        keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, 
        keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, 
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, 
        keyinput31 );
  input N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57,
         N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109,
         N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
         keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10,
         keyinput11, keyinput12, keyinput13, keyinput14, keyinput15,
         keyinput16, keyinput17, keyinput18, keyinput19, keyinput20,
         keyinput21, keyinput22, keyinput23, keyinput24, keyinput25,
         keyinput26, keyinput27, keyinput28, keyinput29, keyinput30,
         keyinput31;
  output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
  wire   n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307;

  XOR2X1 U186 ( .IN1(N125), .IN2(n156), .Q(N755) );
  NOR2X0 U187 ( .IN1(n157), .IN2(n158), .QN(n156) );
  XOR2X1 U188 ( .IN1(N121), .IN2(n159), .Q(N754) );
  NOR2X0 U189 ( .IN1(n160), .IN2(n158), .QN(n159) );
  XOR3X1 U190 ( .IN1(keyinput29), .IN2(N117), .IN3(n161), .Q(N753) );
  OR2X1 U191 ( .IN1(n158), .IN2(n162), .Q(n161) );
  XOR2X1 U192 ( .IN1(N113), .IN2(n163), .Q(N752) );
  NOR2X0 U193 ( .IN1(n164), .IN2(n158), .QN(n163) );
  NAND3X0 U194 ( .IN1(n165), .IN2(n166), .IN3(n167), .QN(n158) );
  XOR3X1 U195 ( .IN1(keyinput28), .IN2(N109), .IN3(n168), .Q(N751) );
  NOR2X0 U196 ( .IN1(n157), .IN2(n169), .QN(n168) );
  XOR2X1 U197 ( .IN1(N105), .IN2(n170), .Q(N750) );
  NOR2X0 U198 ( .IN1(n160), .IN2(n169), .QN(n170) );
  XOR2X1 U199 ( .IN1(N101), .IN2(n171), .Q(N749) );
  NOR2X0 U200 ( .IN1(n162), .IN2(n169), .QN(n171) );
  XOR2X1 U201 ( .IN1(N97), .IN2(n172), .Q(N748) );
  NOR2X0 U202 ( .IN1(n164), .IN2(n169), .QN(n172) );
  NAND3X0 U203 ( .IN1(n165), .IN2(n166), .IN3(n173), .QN(n169) );
  XOR2X1 U204 ( .IN1(N93), .IN2(n174), .Q(N747) );
  NOR2X0 U205 ( .IN1(n157), .IN2(n175), .QN(n174) );
  XOR2X1 U206 ( .IN1(N89), .IN2(n176), .Q(N746) );
  NOR2X0 U207 ( .IN1(n160), .IN2(n175), .QN(n176) );
  XOR3X1 U208 ( .IN1(keyinput27), .IN2(N85), .IN3(n177), .Q(N745) );
  OR2X1 U209 ( .IN1(n175), .IN2(n162), .Q(n177) );
  XOR2X1 U210 ( .IN1(N81), .IN2(n178), .Q(N744) );
  NOR2X0 U211 ( .IN1(n164), .IN2(n175), .QN(n178) );
  NAND3X0 U212 ( .IN1(n167), .IN2(n179), .IN3(n180), .QN(n175) );
  AND3X1 U213 ( .IN1(n181), .IN2(n182), .IN3(n183), .Q(n167) );
  XOR2X1 U214 ( .IN1(N77), .IN2(n184), .Q(N743) );
  NOR2X0 U215 ( .IN1(n157), .IN2(n185), .QN(n184) );
  XOR2X1 U216 ( .IN1(N73), .IN2(n186), .Q(N742) );
  NOR2X0 U217 ( .IN1(n160), .IN2(n185), .QN(n186) );
  XOR2X1 U218 ( .IN1(N69), .IN2(n187), .Q(N741) );
  NOR2X0 U219 ( .IN1(n162), .IN2(n185), .QN(n187) );
  XOR2X1 U220 ( .IN1(N65), .IN2(n188), .Q(N740) );
  NOR2X0 U221 ( .IN1(n164), .IN2(n185), .QN(n188) );
  NAND3X0 U222 ( .IN1(n173), .IN2(n179), .IN3(n180), .QN(n185) );
  AND3X1 U223 ( .IN1(n182), .IN2(n189), .IN3(n190), .Q(n173) );
  XNOR2X1 U224 ( .IN1(n191), .IN2(keyinput23), .Q(n182) );
  NAND3X0 U225 ( .IN1(n192), .IN2(n193), .IN3(n194), .QN(n191) );
  OA222X1 U226 ( .IN1(keyinput21), .IN2(n162), .IN3(n195), .IN4(n157), .IN5(
        keyinput20), .IN6(n196), .Q(n194) );
  OR2X1 U227 ( .IN1(n160), .IN2(keyinput22), .Q(n193) );
  MUX21X1 U228 ( .IN1(n197), .IN2(n198), .S(n164), .Q(n192) );
  OA22X1 U229 ( .IN1(n199), .IN2(n200), .IN3(n201), .IN4(n202), .Q(n198) );
  INVX0 U230 ( .INP(keyinput20), .ZN(n201) );
  AOI22X1 U231 ( .IN1(n162), .IN2(keyinput21), .IN3(keyinput22), .IN4(n160), 
        .QN(n199) );
  AND3X1 U232 ( .IN1(n195), .IN2(n203), .IN3(keyinput20), .Q(n197) );
  NAND3X0 U233 ( .IN1(n157), .IN2(n162), .IN3(n204), .QN(n203) );
  XOR2X1 U234 ( .IN1(keyinput18), .IN2(n205), .Q(n204) );
  AND2X1 U235 ( .IN1(keyinput22), .IN2(keyinput21), .Q(n195) );
  XOR2X1 U236 ( .IN1(N61), .IN2(n206), .Q(N739) );
  NOR2X0 U237 ( .IN1(n190), .IN2(n207), .QN(n206) );
  XOR2X1 U238 ( .IN1(N57), .IN2(n208), .Q(N738) );
  NOR2X0 U239 ( .IN1(n183), .IN2(n207), .QN(n208) );
  XOR2X1 U240 ( .IN1(N53), .IN2(n209), .Q(N737) );
  NOR2X0 U241 ( .IN1(n179), .IN2(n207), .QN(n209) );
  XOR2X1 U242 ( .IN1(N49), .IN2(n210), .Q(N736) );
  NOR2X0 U243 ( .IN1(n166), .IN2(n207), .QN(n210) );
  NAND4X0 U244 ( .IN1(n211), .IN2(n212), .IN3(n200), .IN4(n213), .QN(n207) );
  NOR2X0 U245 ( .IN1(n162), .IN2(n205), .QN(n213) );
  XOR2X1 U246 ( .IN1(keyinput17), .IN2(n164), .Q(n211) );
  XOR2X1 U247 ( .IN1(N45), .IN2(n214), .Q(N735) );
  NOR2X0 U248 ( .IN1(n190), .IN2(n215), .QN(n214) );
  XOR2X1 U249 ( .IN1(N41), .IN2(n216), .Q(N734) );
  NOR2X0 U250 ( .IN1(n183), .IN2(n215), .QN(n216) );
  XOR2X1 U251 ( .IN1(N37), .IN2(n217), .Q(N733) );
  NOR2X0 U252 ( .IN1(n179), .IN2(n215), .QN(n217) );
  XOR2X1 U253 ( .IN1(N33), .IN2(n218), .Q(N732) );
  NOR2X0 U254 ( .IN1(n166), .IN2(n215), .QN(n218) );
  NAND4X0 U255 ( .IN1(n157), .IN2(n212), .IN3(n205), .IN4(n219), .QN(n215) );
  NOR2X0 U256 ( .IN1(n162), .IN2(n220), .QN(n219) );
  XOR2X1 U257 ( .IN1(keyinput16), .IN2(n164), .Q(n220) );
  INVX0 U258 ( .INP(n221), .ZN(n164) );
  XOR3X1 U259 ( .IN1(keyinput26), .IN2(N29), .IN3(n222), .Q(N731) );
  OR2X1 U260 ( .IN1(n223), .IN2(n190), .Q(n222) );
  XOR3X1 U261 ( .IN1(keyinput25), .IN2(N25), .IN3(n224), .Q(N730) );
  NOR2X0 U262 ( .IN1(n183), .IN2(n223), .QN(n224) );
  XOR2X1 U263 ( .IN1(N21), .IN2(n225), .Q(N729) );
  NOR2X0 U264 ( .IN1(n179), .IN2(n223), .QN(n225) );
  XOR2X1 U265 ( .IN1(N17), .IN2(n226), .Q(N728) );
  NOR2X0 U266 ( .IN1(n166), .IN2(n223), .QN(n226) );
  NAND3X0 U267 ( .IN1(n221), .IN2(n212), .IN3(n196), .QN(n223) );
  INVX0 U268 ( .INP(n202), .ZN(n196) );
  NAND3X0 U269 ( .IN1(n200), .IN2(n162), .IN3(n160), .QN(n202) );
  XOR3X1 U270 ( .IN1(keyinput31), .IN2(N13), .IN3(n227), .Q(N727) );
  NAND2X0 U271 ( .IN1(n228), .IN2(n181), .QN(n227) );
  INVX0 U272 ( .INP(n190), .ZN(n181) );
  XOR3X1 U273 ( .IN1(keyinput30), .IN2(N9), .IN3(n229), .Q(N726) );
  NAND2X0 U274 ( .IN1(n228), .IN2(n189), .QN(n229) );
  INVX0 U275 ( .INP(n230), .ZN(n228) );
  XOR2X1 U276 ( .IN1(N5), .IN2(n231), .Q(N725) );
  NOR2X0 U277 ( .IN1(n230), .IN2(n179), .QN(n231) );
  INVX0 U278 ( .INP(n165), .ZN(n179) );
  XOR2X1 U279 ( .IN1(N1), .IN2(n232), .Q(N724) );
  NOR2X0 U280 ( .IN1(n230), .IN2(n166), .QN(n232) );
  XOR2X1 U281 ( .IN1(n233), .IN2(keyinput24), .Q(n230) );
  NAND4X0 U282 ( .IN1(n205), .IN2(n212), .IN3(n221), .IN4(n234), .QN(n233) );
  NOR2X0 U283 ( .IN1(n235), .IN2(n236), .QN(n234) );
  XOR2X1 U284 ( .IN1(keyinput14), .IN2(n162), .Q(n236) );
  XNOR3X1 U285 ( .IN1(n237), .IN2(n238), .IN3(n239), .Q(n162) );
  XOR3X1 U286 ( .IN1(n240), .IN2(n241), .IN3(n242), .Q(n239) );
  NAND2X0 U287 ( .IN1(N134), .IN2(N137), .QN(n241) );
  INVX0 U288 ( .INP(n243), .ZN(n238) );
  XOR2X1 U289 ( .IN1(keyinput15), .IN2(n157), .Q(n235) );
  INVX0 U290 ( .INP(n200), .ZN(n157) );
  XOR3X1 U291 ( .IN1(n244), .IN2(n245), .IN3(n246), .Q(n200) );
  XOR2X1 U292 ( .IN1(n247), .IN2(n248), .Q(n246) );
  INVX0 U293 ( .INP(n240), .ZN(n248) );
  XNOR3X1 U294 ( .IN1(N61), .IN2(N57), .IN3(N49), .Q(n240) );
  XOR3X1 U295 ( .IN1(keyinput10), .IN2(N53), .IN3(n249), .Q(n245) );
  XNOR2X1 U296 ( .IN1(N21), .IN2(n250), .Q(n249) );
  NAND2X0 U297 ( .IN1(N136), .IN2(N137), .QN(n250) );
  XOR2X1 U298 ( .IN1(n251), .IN2(n252), .Q(n244) );
  XOR3X1 U299 ( .IN1(n253), .IN2(n254), .IN3(n255), .Q(n221) );
  XOR3X1 U300 ( .IN1(n247), .IN2(n256), .IN3(n257), .Q(n255) );
  NAND2X0 U301 ( .IN1(N133), .IN2(N137), .QN(n256) );
  XOR3X1 U302 ( .IN1(N25), .IN2(N17), .IN3(n258), .Q(n247) );
  XNOR2X1 U303 ( .IN1(N29), .IN2(keyinput0), .Q(n258) );
  AO21X1 U304 ( .IN1(n190), .IN2(n259), .IN3(n260), .Q(n212) );
  MUX21X1 U305 ( .IN1(n261), .IN2(n262), .S(n263), .Q(n260) );
  NOR3X0 U306 ( .IN1(n264), .IN2(n165), .IN3(n189), .QN(n263) );
  INVX0 U307 ( .INP(n183), .ZN(n189) );
  XOR2X1 U308 ( .IN1(keyinput11), .IN2(n166), .Q(n264) );
  NOR2X0 U309 ( .IN1(n190), .IN2(n261), .QN(n262) );
  AO221X1 U310 ( .IN1(n265), .IN2(n166), .IN3(n266), .IN4(n183), .IN5(n261), 
        .Q(n259) );
  INVX0 U311 ( .INP(keyinput19), .ZN(n261) );
  XOR3X1 U312 ( .IN1(n267), .IN2(n268), .IN3(n269), .Q(n183) );
  XOR3X1 U313 ( .IN1(n270), .IN2(N101), .IN3(n271), .Q(n269) );
  XOR3X1 U314 ( .IN1(N57), .IN2(N41), .IN3(n272), .Q(n271) );
  XOR2X1 U315 ( .IN1(n273), .IN2(N25), .Q(n272) );
  NAND2X0 U316 ( .IN1(N137), .IN2(N131), .QN(n273) );
  XOR3X1 U317 ( .IN1(N77), .IN2(N73), .IN3(n274), .Q(n270) );
  XOR2X1 U318 ( .IN1(keyinput6), .IN2(N9), .Q(n274) );
  XOR3X1 U319 ( .IN1(N69), .IN2(N65), .IN3(n275), .Q(n268) );
  XOR2X1 U320 ( .IN1(keyinput3), .IN2(N97), .Q(n275) );
  XOR2X1 U321 ( .IN1(N109), .IN2(N105), .Q(n267) );
  XOR2X1 U322 ( .IN1(n165), .IN2(n276), .Q(n266) );
  NOR2X0 U323 ( .IN1(keyinput13), .IN2(n166), .QN(n276) );
  INVX0 U324 ( .INP(n180), .ZN(n166) );
  XOR3X1 U325 ( .IN1(n277), .IN2(n278), .IN3(n279), .Q(n180) );
  XNOR2X1 U326 ( .IN1(n257), .IN2(n242), .Q(n279) );
  XNOR3X1 U327 ( .IN1(N85), .IN2(N69), .IN3(N33), .Q(n242) );
  XNOR3X1 U328 ( .IN1(N81), .IN2(N65), .IN3(N1), .Q(n257) );
  XOR3X1 U329 ( .IN1(keyinput9), .IN2(N49), .IN3(n280), .Q(n278) );
  XOR2X1 U330 ( .IN1(n281), .IN2(n282), .Q(n280) );
  NAND2X0 U331 ( .IN1(N129), .IN2(N137), .QN(n282) );
  INVX0 U332 ( .INP(N17), .ZN(n281) );
  XOR2X1 U333 ( .IN1(n251), .IN2(n283), .Q(n277) );
  XOR2X1 U334 ( .IN1(N77), .IN2(N93), .Q(n251) );
  XOR2X1 U335 ( .IN1(n165), .IN2(keyinput12), .Q(n265) );
  XOR3X1 U336 ( .IN1(n237), .IN2(n284), .IN3(n285), .Q(n165) );
  XNOR2X1 U337 ( .IN1(n253), .IN2(n286), .Q(n285) );
  XNOR3X1 U338 ( .IN1(N21), .IN2(N113), .IN3(n287), .Q(n253) );
  XNOR2X1 U339 ( .IN1(N5), .IN2(N97), .Q(n287) );
  XNOR3X1 U340 ( .IN1(keyinput4), .IN2(keyinput3), .IN3(n288), .Q(n284) );
  XOR2X1 U341 ( .IN1(n289), .IN2(n252), .Q(n288) );
  XOR2X1 U342 ( .IN1(N109), .IN2(N125), .Q(n252) );
  NAND2X0 U343 ( .IN1(N130), .IN2(N137), .QN(n289) );
  XNOR3X1 U344 ( .IN1(N117), .IN2(N101), .IN3(n290), .Q(n237) );
  XNOR2X1 U345 ( .IN1(N37), .IN2(N53), .Q(n290) );
  XOR3X1 U346 ( .IN1(n291), .IN2(n292), .IN3(n293), .Q(n190) );
  XOR2X1 U347 ( .IN1(n294), .IN2(n295), .Q(n293) );
  XOR3X1 U348 ( .IN1(N85), .IN2(N81), .IN3(n296), .Q(n295) );
  XOR2X1 U349 ( .IN1(N93), .IN2(N89), .Q(n296) );
  XOR3X1 U350 ( .IN1(N29), .IN2(N13), .IN3(n297), .Q(n294) );
  XNOR2X1 U351 ( .IN1(N45), .IN2(N61), .Q(n297) );
  XOR3X1 U352 ( .IN1(N121), .IN2(N117), .IN3(n298), .Q(n292) );
  XOR2X1 U353 ( .IN1(keyinput4), .IN2(N125), .Q(n298) );
  XOR2X1 U354 ( .IN1(n299), .IN2(n300), .Q(n291) );
  NAND2X0 U355 ( .IN1(N132), .IN2(N137), .QN(n300) );
  INVX0 U356 ( .INP(N113), .ZN(n299) );
  INVX0 U357 ( .INP(n160), .ZN(n205) );
  XOR3X1 U358 ( .IN1(N5), .IN2(N37), .IN3(n301), .Q(n160) );
  XOR3X1 U359 ( .IN1(n302), .IN2(N1), .IN3(n303), .Q(n301) );
  XOR3X1 U360 ( .IN1(n254), .IN2(n304), .IN3(n243), .Q(n303) );
  XOR3X1 U361 ( .IN1(N45), .IN2(N41), .IN3(n305), .Q(n243) );
  XNOR3X1 U362 ( .IN1(keyinput8), .IN2(keyinput2), .IN3(keyinput1), .Q(n305)
         );
  XOR2X1 U363 ( .IN1(n283), .IN2(n286), .Q(n304) );
  XOR2X1 U364 ( .IN1(N105), .IN2(N121), .Q(n286) );
  XOR2X1 U365 ( .IN1(N73), .IN2(N89), .Q(n283) );
  XOR2X1 U366 ( .IN1(N13), .IN2(N9), .Q(n254) );
  XOR3X1 U367 ( .IN1(keyinput7), .IN2(keyinput5), .IN3(n306), .Q(n302) );
  XNOR2X1 U368 ( .IN1(N33), .IN2(n307), .Q(n306) );
  NAND2X0 U369 ( .IN1(N135), .IN2(N137), .QN(n307) );
endmodule

