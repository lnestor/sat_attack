
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436;

  XOR2X1 U281 ( .IN1(n249), .IN2(G32), .Q(G1355) );
  NAND2X0 U282 ( .IN1(n250), .IN2(n251), .QN(n249) );
  XOR2X1 U283 ( .IN1(n252), .IN2(G31), .Q(G1354) );
  NAND2X0 U284 ( .IN1(n250), .IN2(n253), .QN(n252) );
  XOR2X1 U285 ( .IN1(n254), .IN2(G30), .Q(G1353) );
  NAND2X0 U286 ( .IN1(n250), .IN2(n255), .QN(n254) );
  XOR2X1 U287 ( .IN1(n256), .IN2(G29), .Q(G1352) );
  NAND2X0 U288 ( .IN1(n250), .IN2(n257), .QN(n256) );
  AND4X1 U289 ( .IN1(n258), .IN2(n259), .IN3(n260), .IN4(n261), .Q(n250) );
  XOR2X1 U290 ( .IN1(n262), .IN2(n263), .Q(G1351) );
  NOR2X0 U291 ( .IN1(n264), .IN2(n265), .QN(n263) );
  XOR2X1 U292 ( .IN1(n266), .IN2(n267), .Q(G1350) );
  NOR2X0 U293 ( .IN1(n268), .IN2(n265), .QN(n267) );
  XNOR2X1 U294 ( .IN1(G26), .IN2(n269), .Q(G1349) );
  NOR2X0 U295 ( .IN1(n270), .IN2(n265), .QN(n269) );
  XOR2X1 U296 ( .IN1(n271), .IN2(n272), .Q(G1348) );
  NOR2X0 U297 ( .IN1(n273), .IN2(n265), .QN(n272) );
  NAND4X0 U298 ( .IN1(n274), .IN2(n261), .IN3(n260), .IN4(n275), .QN(n265) );
  NOR2X0 U299 ( .IN1(n259), .IN2(n276), .QN(n275) );
  XNOR2X1 U300 ( .IN1(G24), .IN2(n277), .Q(G1347) );
  NOR2X0 U301 ( .IN1(n264), .IN2(n278), .QN(n277) );
  XNOR2X1 U302 ( .IN1(G23), .IN2(n279), .Q(G1346) );
  NOR2X0 U303 ( .IN1(n268), .IN2(n278), .QN(n279) );
  XOR2X1 U304 ( .IN1(n280), .IN2(n281), .Q(G1345) );
  NOR2X0 U305 ( .IN1(n270), .IN2(n278), .QN(n281) );
  XNOR2X1 U306 ( .IN1(G21), .IN2(n282), .Q(G1344) );
  NOR2X0 U307 ( .IN1(n273), .IN2(n278), .QN(n282) );
  NAND4X0 U308 ( .IN1(n276), .IN2(n261), .IN3(n259), .IN4(n283), .QN(n278) );
  NOR2X0 U309 ( .IN1(n260), .IN2(n274), .QN(n283) );
  XOR2X1 U310 ( .IN1(n284), .IN2(G20), .Q(G1343) );
  NAND2X0 U311 ( .IN1(n285), .IN2(n251), .QN(n284) );
  XOR2X1 U312 ( .IN1(n286), .IN2(G19), .Q(G1342) );
  NAND2X0 U313 ( .IN1(n285), .IN2(n253), .QN(n286) );
  XOR2X1 U314 ( .IN1(n287), .IN2(G18), .Q(G1341) );
  NAND2X0 U315 ( .IN1(n285), .IN2(n255), .QN(n287) );
  XOR2X1 U316 ( .IN1(n288), .IN2(G17), .Q(G1340) );
  NAND2X0 U317 ( .IN1(n285), .IN2(n257), .QN(n288) );
  AND4X1 U318 ( .IN1(n289), .IN2(n274), .IN3(n276), .IN4(n261), .Q(n285) );
  NAND2X0 U319 ( .IN1(n290), .IN2(n291), .QN(n261) );
  OR3X1 U320 ( .IN1(n255), .IN2(n292), .IN3(n251), .Q(n291) );
  OR3X1 U321 ( .IN1(n253), .IN2(n293), .IN3(n257), .Q(n290) );
  XOR2X1 U322 ( .IN1(n294), .IN2(G16), .Q(G1339) );
  NAND2X0 U323 ( .IN1(n295), .IN2(n296), .QN(n294) );
  XOR2X1 U324 ( .IN1(n297), .IN2(G15), .Q(G1338) );
  NAND2X0 U325 ( .IN1(n295), .IN2(n298), .QN(n297) );
  XOR2X1 U326 ( .IN1(n299), .IN2(G14), .Q(G1337) );
  NAND2X0 U327 ( .IN1(n295), .IN2(n300), .QN(n299) );
  XOR2X1 U328 ( .IN1(n301), .IN2(G13), .Q(G1336) );
  NAND2X0 U329 ( .IN1(n295), .IN2(n302), .QN(n301) );
  AND4X1 U330 ( .IN1(n293), .IN2(n273), .IN3(n268), .IN4(n303), .Q(n295) );
  NOR2X0 U331 ( .IN1(n270), .IN2(n264), .QN(n293) );
  XNOR2X1 U332 ( .IN1(G12), .IN2(n304), .Q(G1335) );
  NOR2X0 U333 ( .IN1(n274), .IN2(n305), .QN(n304) );
  XNOR2X1 U334 ( .IN1(G11), .IN2(n306), .Q(G1334) );
  NOR2X0 U335 ( .IN1(n259), .IN2(n305), .QN(n306) );
  XNOR2X1 U336 ( .IN1(G10), .IN2(n307), .Q(G1333) );
  NOR2X0 U337 ( .IN1(n276), .IN2(n305), .QN(n307) );
  XNOR2X1 U338 ( .IN1(G9), .IN2(n308), .Q(G1332) );
  NOR2X0 U339 ( .IN1(n260), .IN2(n305), .QN(n308) );
  NAND4X0 U340 ( .IN1(n273), .IN2(n303), .IN3(n264), .IN4(n309), .QN(n305) );
  NOR2X0 U341 ( .IN1(n268), .IN2(n270), .QN(n309) );
  XNOR2X1 U342 ( .IN1(G8), .IN2(n310), .Q(G1331) );
  NOR2X0 U343 ( .IN1(n274), .IN2(n311), .QN(n310) );
  XNOR2X1 U344 ( .IN1(G7), .IN2(n312), .Q(G1330) );
  NOR2X0 U345 ( .IN1(n259), .IN2(n311), .QN(n312) );
  XNOR2X1 U346 ( .IN1(G6), .IN2(n313), .Q(G1329) );
  NOR2X0 U347 ( .IN1(n276), .IN2(n311), .QN(n313) );
  XNOR2X1 U348 ( .IN1(G5), .IN2(n314), .Q(G1328) );
  NOR2X0 U349 ( .IN1(n260), .IN2(n311), .QN(n314) );
  NAND4X0 U350 ( .IN1(n268), .IN2(n303), .IN3(n270), .IN4(n315), .QN(n311) );
  NOR2X0 U351 ( .IN1(n264), .IN2(n273), .QN(n315) );
  XOR2X1 U352 ( .IN1(n316), .IN2(G4), .Q(G1327) );
  NAND2X0 U353 ( .IN1(n317), .IN2(n296), .QN(n316) );
  XOR2X1 U354 ( .IN1(n318), .IN2(G3), .Q(G1326) );
  NAND2X0 U355 ( .IN1(n317), .IN2(n298), .QN(n318) );
  XOR2X1 U356 ( .IN1(n319), .IN2(G2), .Q(G1325) );
  NAND2X0 U357 ( .IN1(n317), .IN2(n300), .QN(n319) );
  XOR2X1 U358 ( .IN1(n320), .IN2(G1), .Q(G1324) );
  NAND2X0 U359 ( .IN1(n317), .IN2(n302), .QN(n320) );
  AND4X1 U360 ( .IN1(n292), .IN2(n264), .IN3(n270), .IN4(n303), .Q(n317) );
  NAND2X0 U361 ( .IN1(n321), .IN2(n322), .QN(n303) );
  OR3X1 U362 ( .IN1(n300), .IN2(n289), .IN3(n296), .Q(n322) );
  NOR2X0 U363 ( .IN1(n260), .IN2(n259), .QN(n289) );
  INVX0 U364 ( .INP(n298), .ZN(n259) );
  INVX0 U365 ( .INP(n302), .ZN(n260) );
  OR3X1 U366 ( .IN1(n302), .IN2(n258), .IN3(n298), .Q(n321) );
  MUX21X1 U367 ( .IN1(n323), .IN2(n324), .S(n325), .Q(n298) );
  XOR3X1 U368 ( .IN1(G15), .IN2(G11), .IN3(n326), .Q(n325) );
  XOR2X1 U369 ( .IN1(G7), .IN2(G3), .Q(n326) );
  NAND2X0 U370 ( .IN1(n327), .IN2(n328), .QN(n324) );
  AND2X1 U371 ( .IN1(n328), .IN2(n327), .Q(n323) );
  NAND3X0 U372 ( .IN1(G35), .IN2(G41), .IN3(n329), .QN(n327) );
  AO21X1 U373 ( .IN1(G35), .IN2(G41), .IN3(n329), .Q(n328) );
  XOR2X1 U374 ( .IN1(n330), .IN2(n331), .Q(n329) );
  NOR2X0 U375 ( .IN1(n276), .IN2(n274), .QN(n258) );
  INVX0 U376 ( .INP(n296), .ZN(n274) );
  MUX21X1 U377 ( .IN1(n332), .IN2(n333), .S(n334), .Q(n296) );
  XOR3X1 U378 ( .IN1(G16), .IN2(G12), .IN3(n335), .Q(n334) );
  XOR2X1 U379 ( .IN1(G8), .IN2(G4), .Q(n335) );
  NAND2X0 U380 ( .IN1(n336), .IN2(n337), .QN(n333) );
  AND2X1 U381 ( .IN1(n337), .IN2(n336), .Q(n332) );
  NAND3X0 U382 ( .IN1(G36), .IN2(G41), .IN3(n338), .QN(n336) );
  AO21X1 U383 ( .IN1(G36), .IN2(G41), .IN3(n338), .Q(n337) );
  XOR2X1 U384 ( .IN1(n339), .IN2(n340), .Q(n338) );
  INVX0 U385 ( .INP(n300), .ZN(n276) );
  MUX21X1 U386 ( .IN1(n341), .IN2(n342), .S(n343), .Q(n300) );
  XOR3X1 U387 ( .IN1(G14), .IN2(G10), .IN3(n344), .Q(n343) );
  XOR2X1 U388 ( .IN1(G6), .IN2(G2), .Q(n344) );
  NAND2X0 U389 ( .IN1(n345), .IN2(n346), .QN(n342) );
  AND2X1 U390 ( .IN1(n346), .IN2(n345), .Q(n341) );
  NAND3X0 U391 ( .IN1(G41), .IN2(n347), .IN3(G34), .QN(n345) );
  AO21X1 U392 ( .IN1(G34), .IN2(G41), .IN3(n347), .Q(n346) );
  XOR2X1 U393 ( .IN1(n340), .IN2(n331), .Q(n347) );
  AND2X1 U394 ( .IN1(n348), .IN2(n349), .Q(n331) );
  XOR2X1 U395 ( .IN1(n350), .IN2(keyinput29), .Q(n349) );
  NAND2X0 U396 ( .IN1(n351), .IN2(n352), .QN(n350) );
  XOR2X1 U397 ( .IN1(n353), .IN2(keyinput30), .Q(n348) );
  NAND2X0 U398 ( .IN1(n352), .IN2(n354), .QN(n353) );
  XNOR2X1 U399 ( .IN1(n355), .IN2(keyinput22), .Q(n352) );
  NAND2X0 U400 ( .IN1(n351), .IN2(n354), .QN(n355) );
  XOR3X1 U401 ( .IN1(keyinput13), .IN2(n262), .IN3(n266), .Q(n354) );
  INVX0 U402 ( .INP(G27), .ZN(n266) );
  INVX0 U403 ( .INP(G28), .ZN(n262) );
  XOR3X1 U404 ( .IN1(keyinput12), .IN2(G26), .IN3(n271), .Q(n351) );
  INVX0 U405 ( .INP(G25), .ZN(n271) );
  AOI21X1 U406 ( .IN1(n356), .IN2(n357), .IN3(n358), .QN(n340) );
  XOR2X1 U407 ( .IN1(keyinput31), .IN2(n359), .Q(n358) );
  AND2X1 U408 ( .IN1(n360), .IN2(n356), .Q(n359) );
  XOR2X1 U409 ( .IN1(n361), .IN2(keyinput23), .Q(n356) );
  NAND2X0 U410 ( .IN1(n360), .IN2(n357), .QN(n361) );
  XOR3X1 U411 ( .IN1(keyinput14), .IN2(G30), .IN3(G29), .Q(n357) );
  XNOR3X1 U412 ( .IN1(keyinput15), .IN2(G32), .IN3(G31), .Q(n360) );
  MUX21X1 U413 ( .IN1(n362), .IN2(n363), .S(n364), .Q(n302) );
  XOR3X1 U414 ( .IN1(G13), .IN2(G1), .IN3(n365), .Q(n364) );
  XOR2X1 U415 ( .IN1(G9), .IN2(G5), .Q(n365) );
  NAND2X0 U416 ( .IN1(n366), .IN2(n367), .QN(n363) );
  AND2X1 U417 ( .IN1(n367), .IN2(n366), .Q(n362) );
  NAND3X0 U418 ( .IN1(G41), .IN2(n368), .IN3(G33), .QN(n366) );
  AO21X1 U419 ( .IN1(G33), .IN2(G41), .IN3(n368), .Q(n367) );
  XOR2X1 U420 ( .IN1(n330), .IN2(n339), .Q(n368) );
  AO21X1 U421 ( .IN1(n369), .IN2(n370), .IN3(n371), .Q(n339) );
  XOR2X1 U422 ( .IN1(n372), .IN2(keyinput21), .Q(n371) );
  OR2X1 U423 ( .IN1(n370), .IN2(n369), .Q(n372) );
  XOR3X1 U424 ( .IN1(keyinput11), .IN2(G24), .IN3(G23), .Q(n370) );
  XOR3X1 U425 ( .IN1(keyinput10), .IN2(n280), .IN3(G21), .Q(n369) );
  INVX0 U426 ( .INP(G22), .ZN(n280) );
  AO21X1 U427 ( .IN1(n373), .IN2(n374), .IN3(n375), .Q(n330) );
  XOR2X1 U428 ( .IN1(keyinput20), .IN2(n376), .Q(n375) );
  NOR2X0 U429 ( .IN1(n373), .IN2(n374), .QN(n376) );
  XNOR3X1 U430 ( .IN1(keyinput9), .IN2(G20), .IN3(G19), .Q(n374) );
  XNOR3X1 U431 ( .IN1(keyinput8), .IN2(G18), .IN3(G17), .Q(n373) );
  INVX0 U432 ( .INP(n255), .ZN(n270) );
  MUX21X1 U433 ( .IN1(n377), .IN2(n378), .S(n379), .Q(n255) );
  XOR3X1 U434 ( .IN1(G22), .IN2(G18), .IN3(n380), .Q(n379) );
  XOR2X1 U435 ( .IN1(G30), .IN2(G26), .Q(n380) );
  NAND2X0 U436 ( .IN1(n381), .IN2(n382), .QN(n378) );
  AND2X1 U437 ( .IN1(n382), .IN2(n381), .Q(n377) );
  NAND3X0 U438 ( .IN1(G38), .IN2(G41), .IN3(n383), .QN(n381) );
  AO21X1 U439 ( .IN1(G38), .IN2(G41), .IN3(n383), .Q(n382) );
  XNOR2X1 U440 ( .IN1(n384), .IN2(n385), .Q(n383) );
  INVX0 U441 ( .INP(n251), .ZN(n264) );
  MUX21X1 U442 ( .IN1(n386), .IN2(n387), .S(n388), .Q(n251) );
  XOR3X1 U443 ( .IN1(G24), .IN2(G20), .IN3(n389), .Q(n388) );
  XOR2X1 U444 ( .IN1(G32), .IN2(G28), .Q(n389) );
  NAND2X0 U445 ( .IN1(n390), .IN2(n391), .QN(n387) );
  AND2X1 U446 ( .IN1(n391), .IN2(n390), .Q(n386) );
  NAND3X0 U447 ( .IN1(G40), .IN2(G41), .IN3(n392), .QN(n390) );
  AO21X1 U448 ( .IN1(G40), .IN2(G41), .IN3(n392), .Q(n391) );
  XOR2X1 U449 ( .IN1(n385), .IN2(n393), .Q(n392) );
  AO21X1 U450 ( .IN1(n394), .IN2(n395), .IN3(n396), .Q(n385) );
  XOR2X1 U451 ( .IN1(n397), .IN2(keyinput19), .Q(n396) );
  OR2X1 U452 ( .IN1(n395), .IN2(n394), .Q(n397) );
  XNOR3X1 U453 ( .IN1(keyinput7), .IN2(G16), .IN3(n398), .Q(n395) );
  INVX0 U454 ( .INP(G15), .ZN(n398) );
  XNOR3X1 U455 ( .IN1(keyinput6), .IN2(G14), .IN3(n399), .Q(n394) );
  INVX0 U456 ( .INP(G13), .ZN(n399) );
  NOR2X0 U457 ( .IN1(n268), .IN2(n273), .QN(n292) );
  INVX0 U458 ( .INP(n257), .ZN(n273) );
  MUX21X1 U459 ( .IN1(n400), .IN2(n401), .S(n402), .Q(n257) );
  XOR3X1 U460 ( .IN1(G21), .IN2(G17), .IN3(n403), .Q(n402) );
  XOR2X1 U461 ( .IN1(G29), .IN2(G25), .Q(n403) );
  NAND2X0 U462 ( .IN1(n404), .IN2(n405), .QN(n401) );
  AND2X1 U463 ( .IN1(n405), .IN2(n404), .Q(n400) );
  NAND3X0 U464 ( .IN1(G41), .IN2(n406), .IN3(G37), .QN(n404) );
  AO21X1 U465 ( .IN1(G37), .IN2(G41), .IN3(n406), .Q(n405) );
  XNOR2X1 U466 ( .IN1(n407), .IN2(n393), .Q(n406) );
  AND2X1 U467 ( .IN1(n408), .IN2(n409), .Q(n393) );
  XOR2X1 U468 ( .IN1(keyinput27), .IN2(n410), .Q(n409) );
  AND2X1 U469 ( .IN1(n411), .IN2(n412), .Q(n410) );
  XOR2X1 U470 ( .IN1(n413), .IN2(keyinput26), .Q(n408) );
  NAND2X0 U471 ( .IN1(n412), .IN2(n414), .QN(n413) );
  XNOR2X1 U472 ( .IN1(n415), .IN2(keyinput17), .Q(n412) );
  NAND2X0 U473 ( .IN1(n414), .IN2(n411), .QN(n415) );
  XOR3X1 U474 ( .IN1(keyinput3), .IN2(G8), .IN3(G7), .Q(n411) );
  XOR3X1 U475 ( .IN1(keyinput2), .IN2(G6), .IN3(G5), .Q(n414) );
  INVX0 U476 ( .INP(n253), .ZN(n268) );
  MUX21X1 U477 ( .IN1(n416), .IN2(n417), .S(n418), .Q(n253) );
  XOR3X1 U478 ( .IN1(G23), .IN2(G19), .IN3(n419), .Q(n418) );
  XOR2X1 U479 ( .IN1(G31), .IN2(G27), .Q(n419) );
  NAND2X0 U480 ( .IN1(n420), .IN2(n421), .QN(n417) );
  AND2X1 U481 ( .IN1(n421), .IN2(n420), .Q(n416) );
  NAND3X0 U482 ( .IN1(G39), .IN2(n422), .IN3(G41), .QN(n420) );
  AO21X1 U483 ( .IN1(G41), .IN2(G39), .IN3(n422), .Q(n421) );
  XOR2X1 U484 ( .IN1(n407), .IN2(n384), .Q(n422) );
  AO21X1 U485 ( .IN1(n423), .IN2(n424), .IN3(n425), .Q(n384) );
  XOR2X1 U486 ( .IN1(n426), .IN2(keyinput28), .Q(n425) );
  NAND2X0 U487 ( .IN1(n423), .IN2(n427), .QN(n426) );
  XOR2X1 U488 ( .IN1(n428), .IN2(keyinput18), .Q(n423) );
  NAND2X0 U489 ( .IN1(n427), .IN2(n424), .QN(n428) );
  XOR3X1 U490 ( .IN1(keyinput5), .IN2(G12), .IN3(G11), .Q(n424) );
  XNOR3X1 U491 ( .IN1(keyinput4), .IN2(G9), .IN3(G10), .Q(n427) );
  NAND2X0 U492 ( .IN1(n429), .IN2(n430), .QN(n407) );
  XOR2X1 U493 ( .IN1(n431), .IN2(keyinput25), .Q(n430) );
  NAND2X0 U494 ( .IN1(n432), .IN2(n433), .QN(n431) );
  XOR2X1 U495 ( .IN1(n434), .IN2(keyinput24), .Q(n429) );
  NAND2X0 U496 ( .IN1(n432), .IN2(n435), .QN(n434) );
  XNOR2X1 U497 ( .IN1(n436), .IN2(keyinput16), .Q(n432) );
  NAND2X0 U498 ( .IN1(n435), .IN2(n433), .QN(n436) );
  XOR3X1 U499 ( .IN1(keyinput1), .IN2(G4), .IN3(G3), .Q(n433) );
  XOR3X1 U500 ( .IN1(keyinput0), .IN2(G2), .IN3(G1), .Q(n435) );
endmodule

