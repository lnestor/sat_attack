
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133;

  XOR2X1 U594 ( .IN1(keyinput255), .IN2(n573), .Q(G1351) );
  NOR2X0 U595 ( .IN1(n574), .IN2(n575), .QN(n573) );
  XOR2X1 U596 ( .IN1(n576), .IN2(keyinput220), .Q(n575) );
  NAND3X0 U597 ( .IN1(n577), .IN2(n578), .IN3(n579), .QN(n576) );
  OA21X1 U598 ( .IN1(n580), .IN2(n581), .IN3(G28), .Q(n574) );
  XNOR2X1 U599 ( .IN1(n582), .IN2(keyinput252), .Q(G1346) );
  NAND2X0 U600 ( .IN1(n583), .IN2(n584), .QN(n582) );
  NAND3X0 U601 ( .IN1(n585), .IN2(n586), .IN3(n587), .QN(n584) );
  XOR2X1 U602 ( .IN1(keyinput217), .IN2(n588), .Q(n583) );
  AND2X1 U603 ( .IN1(n587), .IN2(G23), .Q(n588) );
  XNOR2X1 U604 ( .IN1(n589), .IN2(keyinput196), .Q(n587) );
  NAND3X0 U605 ( .IN1(n585), .IN2(n586), .IN3(G23), .QN(n589) );
  XNOR3X1 U606 ( .IN1(keyinput251), .IN2(keyinput234), .IN3(n590), .Q(G1345)
         );
  NOR2X0 U607 ( .IN1(n591), .IN2(n592), .QN(n590) );
  XOR2X1 U608 ( .IN1(n593), .IN2(keyinput216), .Q(n592) );
  NAND3X0 U609 ( .IN1(n594), .IN2(n595), .IN3(n585), .QN(n593) );
  AOI21X1 U610 ( .IN1(n594), .IN2(n585), .IN3(n595), .QN(n591) );
  XOR3X1 U611 ( .IN1(keyinput250), .IN2(keyinput232), .IN3(n596), .Q(G1343) );
  NAND2X0 U612 ( .IN1(n597), .IN2(n598), .QN(n596) );
  XOR2X1 U613 ( .IN1(keyinput215), .IN2(n599), .Q(n598) );
  NOR2X0 U614 ( .IN1(G20), .IN2(n600), .QN(n599) );
  XOR2X1 U615 ( .IN1(n601), .IN2(keyinput214), .Q(n597) );
  NAND2X0 U616 ( .IN1(G20), .IN2(n600), .QN(n601) );
  NAND2X0 U617 ( .IN1(n602), .IN2(n577), .QN(n600) );
  XOR3X1 U618 ( .IN1(keyinput241), .IN2(keyinput226), .IN3(n603), .Q(G1331) );
  OA21X1 U619 ( .IN1(n604), .IN2(n605), .IN3(n606), .Q(n603) );
  XOR2X1 U620 ( .IN1(keyinput205), .IN2(n607), .Q(n606) );
  NOR2X0 U621 ( .IN1(n604), .IN2(n608), .QN(n607) );
  XOR2X1 U622 ( .IN1(n609), .IN2(keyinput185), .Q(n604) );
  OR2X1 U623 ( .IN1(n608), .IN2(n605), .Q(n609) );
  XNOR2X1 U624 ( .IN1(n610), .IN2(keyinput174), .Q(n608) );
  NAND2X0 U625 ( .IN1(n611), .IN2(n612), .QN(n610) );
  XNOR3X1 U626 ( .IN1(n613), .IN2(G5), .IN3(n614), .Q(G1328) );
  NAND2X0 U627 ( .IN1(n611), .IN2(n615), .QN(n614) );
  XOR3X1 U628 ( .IN1(keyinput238), .IN2(keyinput225), .IN3(keyinput172), .Q(
        n613) );
  XNOR2X1 U629 ( .IN1(keyinput235), .IN2(n616), .Q(G1355) );
  OA21X1 U630 ( .IN1(n617), .IN2(n618), .IN3(n619), .Q(n616) );
  XOR2X1 U631 ( .IN1(keyinput224), .IN2(n620), .Q(n619) );
  NOR2X0 U632 ( .IN1(n621), .IN2(n618), .QN(n620) );
  XNOR2X1 U633 ( .IN1(n622), .IN2(keyinput201), .Q(n618) );
  OR2X1 U634 ( .IN1(n621), .IN2(n617), .Q(n622) );
  XNOR2X1 U635 ( .IN1(n623), .IN2(keyinput181), .Q(n621) );
  NAND2X0 U636 ( .IN1(n624), .IN2(n577), .QN(n623) );
  OAI21X1 U637 ( .IN1(n625), .IN2(G31), .IN3(n626), .QN(G1354) );
  XNOR2X1 U638 ( .IN1(n627), .IN2(keyinput200), .Q(n626) );
  NAND2X0 U639 ( .IN1(G31), .IN2(n625), .QN(n627) );
  XNOR2X1 U640 ( .IN1(n628), .IN2(keyinput180), .Q(n625) );
  NAND2X0 U641 ( .IN1(n624), .IN2(n586), .QN(n628) );
  NOR2X0 U642 ( .IN1(n629), .IN2(n630), .QN(G1353) );
  XOR2X1 U643 ( .IN1(keyinput223), .IN2(n631), .Q(n630) );
  NOR2X0 U644 ( .IN1(G30), .IN2(n632), .QN(n631) );
  XOR2X1 U645 ( .IN1(n633), .IN2(keyinput222), .Q(n629) );
  NAND2X0 U646 ( .IN1(G30), .IN2(n632), .QN(n633) );
  NAND2X0 U647 ( .IN1(n624), .IN2(n594), .QN(n632) );
  OA21X1 U648 ( .IN1(n634), .IN2(n635), .IN3(n636), .Q(G1352) );
  XOR2X1 U649 ( .IN1(keyinput221), .IN2(n637), .Q(n636) );
  NOR2X0 U650 ( .IN1(n634), .IN2(n638), .QN(n637) );
  XOR2X1 U651 ( .IN1(n639), .IN2(keyinput199), .Q(n634) );
  OR2X1 U652 ( .IN1(n638), .IN2(n635), .Q(n639) );
  NAND2X0 U653 ( .IN1(n624), .IN2(n640), .QN(n638) );
  XOR2X1 U654 ( .IN1(n641), .IN2(keyinput169), .Q(n624) );
  NAND3X0 U655 ( .IN1(n642), .IN2(n643), .IN3(n644), .QN(n641) );
  OA21X1 U656 ( .IN1(n645), .IN2(n646), .IN3(n647), .Q(G1349) );
  XOR2X1 U657 ( .IN1(n648), .IN2(keyinput218), .Q(n647) );
  NAND3X0 U658 ( .IN1(n594), .IN2(n646), .IN3(n579), .QN(n648) );
  NOR2X0 U659 ( .IN1(n649), .IN2(n581), .QN(n645) );
  AO21X1 U660 ( .IN1(n650), .IN2(n651), .IN3(n652), .Q(G1348) );
  XOR2X1 U661 ( .IN1(n653), .IN2(keyinput198), .Q(n652) );
  OR2X1 U662 ( .IN1(n650), .IN2(n651), .Q(n653) );
  XNOR2X1 U663 ( .IN1(n654), .IN2(keyinput179), .Q(n650) );
  NAND2X0 U664 ( .IN1(n579), .IN2(n640), .QN(n654) );
  INVX0 U665 ( .INP(n581), .ZN(n579) );
  NOR2X0 U666 ( .IN1(n655), .IN2(n656), .QN(G1338) );
  XOR2X1 U667 ( .IN1(keyinput210), .IN2(n657), .Q(n656) );
  AND2X1 U668 ( .IN1(n658), .IN2(G15), .Q(n657) );
  XOR2X1 U669 ( .IN1(n659), .IN2(keyinput211), .Q(n655) );
  NAND2X0 U670 ( .IN1(n660), .IN2(n658), .QN(n659) );
  XNOR2X1 U671 ( .IN1(n661), .IN2(keyinput191), .Q(n658) );
  NAND2X0 U672 ( .IN1(n660), .IN2(G15), .QN(n661) );
  AND2X1 U673 ( .IN1(n662), .IN2(n663), .Q(n660) );
  OA22X1 U674 ( .IN1(n664), .IN2(n665), .IN3(n664), .IN4(n666), .Q(G1335) );
  XOR2X1 U675 ( .IN1(n667), .IN2(keyinput188), .Q(n664) );
  OR2X1 U676 ( .IN1(n665), .IN2(n666), .Q(n667) );
  NAND2X0 U677 ( .IN1(n612), .IN2(n668), .QN(n665) );
  XOR2X1 U678 ( .IN1(n669), .IN2(n670), .Q(G1334) );
  AND2X1 U679 ( .IN1(n663), .IN2(n668), .Q(n670) );
  AO21X1 U680 ( .IN1(n671), .IN2(n672), .IN3(n673), .Q(G1325) );
  XOR2X1 U681 ( .IN1(keyinput182), .IN2(n674), .Q(n673) );
  NOR2X0 U682 ( .IN1(n671), .IN2(n672), .QN(n674) );
  INVX0 U683 ( .INP(G2), .ZN(n672) );
  XOR2X1 U684 ( .IN1(n675), .IN2(keyinput170), .Q(n671) );
  NAND2X0 U685 ( .IN1(n676), .IN2(n642), .QN(n675) );
  NOR2X0 U686 ( .IN1(n677), .IN2(n678), .QN(G1324) );
  XOR2X1 U687 ( .IN1(n679), .IN2(keyinput203), .Q(n678) );
  OR2X1 U688 ( .IN1(n680), .IN2(G1), .Q(n679) );
  XOR2X1 U689 ( .IN1(n681), .IN2(keyinput202), .Q(n677) );
  NAND2X0 U690 ( .IN1(G1), .IN2(n680), .QN(n681) );
  NAND2X0 U691 ( .IN1(n676), .IN2(n615), .QN(n680) );
  XOR2X1 U692 ( .IN1(keyinput233), .IN2(n682), .Q(G1344) );
  OA21X1 U693 ( .IN1(G21), .IN2(n683), .IN3(n684), .Q(n682) );
  XOR2X1 U694 ( .IN1(keyinput195), .IN2(n685), .Q(n684) );
  AND2X1 U695 ( .IN1(n683), .IN2(G21), .Q(n685) );
  XNOR2X1 U696 ( .IN1(n686), .IN2(keyinput177), .Q(n683) );
  NAND2X0 U697 ( .IN1(n585), .IN2(n640), .QN(n686) );
  XOR2X1 U698 ( .IN1(keyinput254), .IN2(n687), .Q(G1350) );
  NOR2X0 U699 ( .IN1(n688), .IN2(n689), .QN(n687) );
  XOR2X1 U700 ( .IN1(n690), .IN2(keyinput219), .Q(n689) );
  OR3X1 U701 ( .IN1(n691), .IN2(G27), .IN3(n581), .Q(n690) );
  OA21X1 U702 ( .IN1(n691), .IN2(n581), .IN3(G27), .Q(n688) );
  NAND4X0 U703 ( .IN1(n663), .IN2(n692), .IN3(n693), .IN4(n694), .QN(n581) );
  NOR2X0 U704 ( .IN1(n695), .IN2(n696), .QN(n694) );
  XOR2X1 U705 ( .IN1(n615), .IN2(keyinput157), .Q(n695) );
  XOR2X1 U706 ( .IN1(keyinput253), .IN2(n697), .Q(G1347) );
  OA21X1 U707 ( .IN1(G24), .IN2(n698), .IN3(n699), .Q(n697) );
  XOR2X1 U708 ( .IN1(n700), .IN2(keyinput197), .Q(n699) );
  NAND2X0 U709 ( .IN1(G24), .IN2(n698), .QN(n700) );
  XNOR2X1 U710 ( .IN1(n701), .IN2(keyinput178), .Q(n698) );
  NAND2X0 U711 ( .IN1(n577), .IN2(n585), .QN(n701) );
  XNOR2X1 U712 ( .IN1(n702), .IN2(keyinput168), .Q(n585) );
  NAND3X0 U713 ( .IN1(n696), .IN2(n615), .IN3(n644), .QN(n702) );
  AND3X1 U714 ( .IN1(n612), .IN2(n692), .IN3(n703), .Q(n644) );
  XNOR3X1 U715 ( .IN1(keyinput249), .IN2(keyinput231), .IN3(n704), .Q(G1342)
         );
  OA22X1 U716 ( .IN1(n705), .IN2(n706), .IN3(n707), .IN4(n706), .Q(n704) );
  XNOR2X1 U717 ( .IN1(n708), .IN2(keyinput194), .Q(n706) );
  OR2X1 U718 ( .IN1(n705), .IN2(n707), .Q(n708) );
  NAND2X0 U719 ( .IN1(n602), .IN2(n586), .QN(n705) );
  XNOR2X1 U720 ( .IN1(keyinput248), .IN2(n709), .Q(G1341) );
  AOI21X1 U721 ( .IN1(n710), .IN2(n711), .IN3(n712), .QN(n709) );
  XNOR2X1 U722 ( .IN1(n713), .IN2(keyinput213), .Q(n712) );
  NAND2X0 U723 ( .IN1(n711), .IN2(G18), .QN(n713) );
  XOR2X1 U724 ( .IN1(n714), .IN2(keyinput193), .Q(n711) );
  NAND2X0 U725 ( .IN1(n710), .IN2(G18), .QN(n714) );
  XOR2X1 U726 ( .IN1(n715), .IN2(keyinput176), .Q(n710) );
  NAND2X0 U727 ( .IN1(n602), .IN2(n594), .QN(n715) );
  XOR2X1 U728 ( .IN1(keyinput247), .IN2(n716), .Q(G1340) );
  OA21X1 U729 ( .IN1(G17), .IN2(n717), .IN3(n718), .Q(n716) );
  XOR2X1 U730 ( .IN1(n719), .IN2(keyinput212), .Q(n718) );
  NAND2X0 U731 ( .IN1(G17), .IN2(n717), .QN(n719) );
  XNOR2X1 U732 ( .IN1(n720), .IN2(keyinput175), .Q(n717) );
  NAND2X0 U733 ( .IN1(n602), .IN2(n640), .QN(n720) );
  AND4X1 U734 ( .IN1(n615), .IN2(n692), .IN3(n696), .IN4(n721), .Q(n602) );
  NOR2X0 U735 ( .IN1(n703), .IN2(n612), .QN(n721) );
  NAND4X0 U736 ( .IN1(n722), .IN2(n723), .IN3(n724), .IN4(n725), .QN(n692) );
  XNOR2X1 U737 ( .IN1(n726), .IN2(keyinput160), .Q(n725) );
  NAND4X0 U738 ( .IN1(n691), .IN2(n577), .IN3(n727), .IN4(n728), .QN(n726) );
  XOR2X1 U739 ( .IN1(keyinput151), .IN2(n729), .Q(n728) );
  XOR2X1 U740 ( .IN1(keyinput152), .IN2(n594), .Q(n727) );
  XNOR2X1 U741 ( .IN1(n730), .IN2(keyinput162), .Q(n724) );
  NAND4X0 U742 ( .IN1(n731), .IN2(n691), .IN3(n732), .IN4(n594), .QN(n730) );
  XOR2X1 U743 ( .IN1(keyinput153), .IN2(n729), .Q(n732) );
  XOR2X1 U744 ( .IN1(n577), .IN2(keyinput154), .Q(n731) );
  XNOR2X1 U745 ( .IN1(n733), .IN2(keyinput163), .Q(n723) );
  NAND4X0 U746 ( .IN1(n734), .IN2(n735), .IN3(n580), .IN4(n640), .QN(n733) );
  INVX0 U747 ( .INP(n577), .ZN(n580) );
  XOR2X1 U748 ( .IN1(keyinput155), .IN2(n594), .Q(n735) );
  XOR2X1 U749 ( .IN1(n691), .IN2(keyinput156), .Q(n734) );
  XOR2X1 U750 ( .IN1(n736), .IN2(keyinput161), .Q(n722) );
  NAND2X0 U751 ( .IN1(n737), .IN2(n729), .QN(n736) );
  XNOR3X1 U752 ( .IN1(keyinput246), .IN2(keyinput230), .IN3(n738), .Q(G1339)
         );
  AOI21X1 U753 ( .IN1(n739), .IN2(G16), .IN3(n740), .QN(n738) );
  AND3X1 U754 ( .IN1(n612), .IN2(n739), .IN3(n662), .Q(n740) );
  XNOR2X1 U755 ( .IN1(n741), .IN2(keyinput192), .Q(n739) );
  NAND3X0 U756 ( .IN1(n612), .IN2(G16), .IN3(n662), .QN(n741) );
  XNOR3X1 U757 ( .IN1(keyinput245), .IN2(keyinput229), .IN3(n742), .Q(G1337)
         );
  AOI21X1 U758 ( .IN1(G14), .IN2(n743), .IN3(n744), .QN(n742) );
  XNOR2X1 U759 ( .IN1(n745), .IN2(keyinput209), .Q(n744) );
  NAND2X0 U760 ( .IN1(n743), .IN2(n746), .QN(n745) );
  XOR2X1 U761 ( .IN1(n747), .IN2(keyinput190), .Q(n743) );
  NAND2X0 U762 ( .IN1(n746), .IN2(G14), .QN(n747) );
  AND2X1 U763 ( .IN1(n662), .IN2(n642), .Q(n746) );
  XNOR2X1 U764 ( .IN1(keyinput244), .IN2(n748), .Q(G1336) );
  OA21X1 U765 ( .IN1(n749), .IN2(n750), .IN3(n751), .Q(n748) );
  XOR2X1 U766 ( .IN1(keyinput208), .IN2(n752), .Q(n751) );
  NOR2X0 U767 ( .IN1(n749), .IN2(n753), .QN(n752) );
  XOR2X1 U768 ( .IN1(n754), .IN2(keyinput189), .Q(n749) );
  OR2X1 U769 ( .IN1(n753), .IN2(n750), .Q(n754) );
  INVX0 U770 ( .INP(G13), .ZN(n750) );
  NAND2X0 U771 ( .IN1(n662), .IN2(n615), .QN(n753) );
  XOR2X1 U772 ( .IN1(n755), .IN2(keyinput167), .Q(n662) );
  NAND3X0 U773 ( .IN1(n691), .IN2(n577), .IN3(n756), .QN(n755) );
  XOR3X1 U774 ( .IN1(keyinput243), .IN2(keyinput228), .IN3(n757), .Q(G1333) );
  OA21X1 U775 ( .IN1(n758), .IN2(n759), .IN3(n760), .Q(n757) );
  XOR2X1 U776 ( .IN1(keyinput207), .IN2(n761), .Q(n760) );
  NOR2X0 U777 ( .IN1(n762), .IN2(n759), .QN(n761) );
  XNOR2X1 U778 ( .IN1(n763), .IN2(keyinput187), .Q(n759) );
  OR2X1 U779 ( .IN1(n762), .IN2(n758), .Q(n763) );
  NAND2X0 U780 ( .IN1(n642), .IN2(n668), .QN(n762) );
  XOR3X1 U781 ( .IN1(keyinput242), .IN2(keyinput227), .IN3(n764), .Q(G1332) );
  NAND2X0 U782 ( .IN1(n765), .IN2(n766), .QN(n764) );
  NAND3X0 U783 ( .IN1(n668), .IN2(n615), .IN3(n767), .QN(n766) );
  XOR2X1 U784 ( .IN1(keyinput206), .IN2(n768), .Q(n765) );
  AND2X1 U785 ( .IN1(n767), .IN2(G9), .Q(n768) );
  XNOR2X1 U786 ( .IN1(n769), .IN2(keyinput186), .Q(n767) );
  NAND3X0 U787 ( .IN1(n668), .IN2(n615), .IN3(G9), .QN(n769) );
  XNOR2X1 U788 ( .IN1(n770), .IN2(keyinput166), .Q(n668) );
  NAND3X0 U789 ( .IN1(n756), .IN2(n586), .IN3(n771), .QN(n770) );
  XOR2X1 U790 ( .IN1(n577), .IN2(keyinput150), .Q(n771) );
  AND3X1 U791 ( .IN1(n729), .IN2(n594), .IN3(n772), .Q(n756) );
  INVX0 U792 ( .INP(n640), .ZN(n729) );
  XNOR2X1 U793 ( .IN1(keyinput240), .IN2(n773), .Q(G1330) );
  OA21X1 U794 ( .IN1(n774), .IN2(n775), .IN3(n776), .Q(n773) );
  XOR2X1 U795 ( .IN1(n777), .IN2(keyinput204), .Q(n776) );
  NAND2X0 U796 ( .IN1(n778), .IN2(n779), .QN(n777) );
  INVX0 U797 ( .INP(n774), .ZN(n779) );
  XOR2X1 U798 ( .IN1(n780), .IN2(keyinput184), .Q(n774) );
  NAND2X0 U799 ( .IN1(n778), .IN2(G7), .QN(n780) );
  AND2X1 U800 ( .IN1(n611), .IN2(n663), .Q(n778) );
  XOR2X1 U801 ( .IN1(keyinput239), .IN2(n781), .Q(G1329) );
  OA21X1 U802 ( .IN1(G6), .IN2(n782), .IN3(n783), .Q(n781) );
  XOR2X1 U803 ( .IN1(keyinput183), .IN2(n784), .Q(n783) );
  AND2X1 U804 ( .IN1(G6), .IN2(n782), .Q(n784) );
  XOR2X1 U805 ( .IN1(n785), .IN2(keyinput173), .Q(n782) );
  NAND2X0 U806 ( .IN1(n611), .IN2(n642), .QN(n785) );
  AND4X1 U807 ( .IN1(n786), .IN2(n640), .IN3(n691), .IN4(n787), .Q(n611) );
  AND2X1 U808 ( .IN1(n577), .IN2(n772), .Q(n787) );
  XOR2X1 U809 ( .IN1(keyinput149), .IN2(n594), .Q(n786) );
  XOR3X1 U810 ( .IN1(keyinput237), .IN2(n788), .IN3(n789), .Q(G1327) );
  NAND2X0 U811 ( .IN1(n676), .IN2(n612), .QN(n789) );
  XOR3X1 U812 ( .IN1(G3), .IN2(n790), .IN3(n791), .Q(G1326) );
  NAND2X0 U813 ( .IN1(n676), .IN2(n663), .QN(n791) );
  INVX0 U814 ( .INP(n703), .ZN(n663) );
  XOR2X1 U815 ( .IN1(n792), .IN2(keyinput165), .Q(n676) );
  NAND4X0 U816 ( .IN1(n772), .IN2(n737), .IN3(n586), .IN4(n640), .QN(n792) );
  AO21X1 U817 ( .IN1(n793), .IN2(n794), .IN3(n795), .Q(n640) );
  XOR2X1 U818 ( .IN1(n796), .IN2(keyinput136), .Q(n795) );
  NAND2X0 U819 ( .IN1(n793), .IN2(n797), .QN(n796) );
  XNOR2X1 U820 ( .IN1(n798), .IN2(keyinput129), .Q(n793) );
  NAND2X0 U821 ( .IN1(n794), .IN2(n797), .QN(n798) );
  OAI21X1 U822 ( .IN1(n799), .IN2(keyinput118), .IN3(n800), .QN(n797) );
  XNOR2X1 U823 ( .IN1(n801), .IN2(n802), .Q(n800) );
  NAND2X0 U824 ( .IN1(keyinput118), .IN2(n799), .QN(n802) );
  NAND2X0 U825 ( .IN1(G37), .IN2(G41), .QN(n801) );
  AO21X1 U826 ( .IN1(n803), .IN2(n804), .IN3(n805), .Q(n799) );
  XOR2X1 U827 ( .IN1(n806), .IN2(keyinput99), .Q(n805) );
  OR2X1 U828 ( .IN1(n804), .IN2(n803), .Q(n806) );
  XNOR3X1 U829 ( .IN1(n807), .IN2(n808), .IN3(n809), .Q(n794) );
  XNOR2X1 U830 ( .IN1(keyinput92), .IN2(keyinput61), .Q(n809) );
  NOR2X0 U831 ( .IN1(n810), .IN2(n811), .QN(n808) );
  XOR2X1 U832 ( .IN1(keyinput38), .IN2(n812), .Q(n811) );
  NOR2X0 U833 ( .IN1(n813), .IN2(n814), .QN(n812) );
  XOR2X1 U834 ( .IN1(keyinput37), .IN2(n815), .Q(n810) );
  NOR2X0 U835 ( .IN1(n813), .IN2(n816), .QN(n815) );
  INVX0 U836 ( .INP(G17), .ZN(n816) );
  XOR2X1 U837 ( .IN1(n817), .IN2(keyinput13), .Q(n813) );
  NAND2X0 U838 ( .IN1(G21), .IN2(G17), .QN(n817) );
  OA21X1 U839 ( .IN1(n818), .IN2(n635), .IN3(n819), .Q(n807) );
  XOR2X1 U840 ( .IN1(keyinput39), .IN2(n820), .Q(n819) );
  NOR2X0 U841 ( .IN1(n818), .IN2(n651), .QN(n820) );
  XOR2X1 U842 ( .IN1(n821), .IN2(keyinput14), .Q(n818) );
  NAND2X0 U843 ( .IN1(G29), .IN2(G25), .QN(n821) );
  INVX0 U844 ( .INP(n691), .ZN(n586) );
  XNOR3X1 U845 ( .IN1(keyinput94), .IN2(n822), .IN3(n823), .Q(n691) );
  OA21X1 U846 ( .IN1(n824), .IN2(n825), .IN3(n826), .Q(n823) );
  XOR2X1 U847 ( .IN1(n827), .IN2(keyinput81), .Q(n826) );
  NAND2X0 U848 ( .IN1(n828), .IN2(n829), .QN(n827) );
  INVX0 U849 ( .INP(n828), .ZN(n825) );
  XOR2X1 U850 ( .IN1(n830), .IN2(keyinput69), .Q(n828) );
  NAND2X0 U851 ( .IN1(n831), .IN2(n829), .QN(n830) );
  AO21X1 U852 ( .IN1(n832), .IN2(G31), .IN3(n833), .Q(n829) );
  XOR2X1 U853 ( .IN1(keyinput42), .IN2(n834), .Q(n833) );
  AND2X1 U854 ( .IN1(G27), .IN2(n832), .Q(n834) );
  XOR2X1 U855 ( .IN1(n835), .IN2(keyinput17), .Q(n832) );
  NAND2X0 U856 ( .IN1(G31), .IN2(G27), .QN(n835) );
  INVX0 U857 ( .INP(n824), .ZN(n831) );
  AO21X1 U858 ( .IN1(n707), .IN2(n836), .IN3(n837), .Q(n824) );
  XOR2X1 U859 ( .IN1(keyinput16), .IN2(n838), .Q(n837) );
  NOR2X0 U860 ( .IN1(n707), .IN2(n836), .QN(n838) );
  OA21X1 U861 ( .IN1(n839), .IN2(n840), .IN3(n841), .Q(n822) );
  XOR2X1 U862 ( .IN1(keyinput121), .IN2(n842), .Q(n841) );
  NOR2X0 U863 ( .IN1(n840), .IN2(n843), .QN(n842) );
  XOR2X1 U864 ( .IN1(n844), .IN2(keyinput114), .Q(n840) );
  OR2X1 U865 ( .IN1(n843), .IN2(n839), .Q(n844) );
  XNOR2X1 U866 ( .IN1(n845), .IN2(keyinput2), .Q(n843) );
  NAND2X0 U867 ( .IN1(G39), .IN2(G41), .QN(n845) );
  XNOR3X1 U868 ( .IN1(keyinput108), .IN2(n804), .IN3(n846), .Q(n839) );
  XOR2X1 U869 ( .IN1(keyinput83), .IN2(n847), .Q(n804) );
  OA21X1 U870 ( .IN1(n848), .IN2(n849), .IN3(n850), .Q(n847) );
  XOR2X1 U871 ( .IN1(keyinput70), .IN2(n851), .Q(n850) );
  NOR2X0 U872 ( .IN1(n848), .IN2(n852), .QN(n851) );
  NOR2X0 U873 ( .IN1(n849), .IN2(n852), .QN(n848) );
  AOI21X1 U874 ( .IN1(n853), .IN2(G1), .IN3(n854), .QN(n852) );
  XOR2X1 U875 ( .IN1(n855), .IN2(keyinput19), .Q(n854) );
  NAND2X0 U876 ( .IN1(n853), .IN2(G2), .QN(n855) );
  XOR2X1 U877 ( .IN1(n856), .IN2(keyinput3), .Q(n853) );
  NAND2X0 U878 ( .IN1(G2), .IN2(G1), .QN(n856) );
  XNOR2X1 U879 ( .IN1(keyinput46), .IN2(n857), .Q(n849) );
  OA21X1 U880 ( .IN1(G3), .IN2(n788), .IN3(n858), .Q(n857) );
  XOR2X1 U881 ( .IN1(keyinput20), .IN2(n859), .Q(n858) );
  NOR2X0 U882 ( .IN1(G4), .IN2(n860), .QN(n859) );
  INVX0 U883 ( .INP(G4), .ZN(n788) );
  NOR2X0 U884 ( .IN1(n594), .IN2(n577), .QN(n737) );
  XOR3X1 U885 ( .IN1(n861), .IN2(n862), .IN3(n863), .Q(n577) );
  XNOR3X1 U886 ( .IN1(keyinput95), .IN2(keyinput142), .IN3(keyinput126), .Q(
        n863) );
  OA21X1 U887 ( .IN1(n864), .IN2(n865), .IN3(n866), .Q(n862) );
  XOR2X1 U888 ( .IN1(n867), .IN2(n868), .Q(n866) );
  AND2X1 U889 ( .IN1(n865), .IN2(n864), .Q(n868) );
  NAND2X0 U890 ( .IN1(G41), .IN2(G40), .QN(n867) );
  INVX0 U891 ( .INP(keyinput122), .ZN(n865) );
  XOR2X1 U892 ( .IN1(keyinput109), .IN2(n869), .Q(n864) );
  OA21X1 U893 ( .IN1(n870), .IN2(n871), .IN3(n872), .Q(n869) );
  XOR2X1 U894 ( .IN1(n873), .IN2(keyinput101), .Q(n872) );
  NAND2X0 U895 ( .IN1(n870), .IN2(n871), .QN(n873) );
  INVX0 U896 ( .INP(n803), .ZN(n871) );
  XNOR3X1 U897 ( .IN1(n874), .IN2(n875), .IN3(G5), .Q(n803) );
  XOR3X1 U898 ( .IN1(keyinput84), .IN2(keyinput47), .IN3(G6), .Q(n875) );
  OA21X1 U899 ( .IN1(G8), .IN2(n775), .IN3(n876), .Q(n874) );
  XOR2X1 U900 ( .IN1(n877), .IN2(keyinput21), .Q(n876) );
  NAND2X0 U901 ( .IN1(G8), .IN2(n775), .QN(n877) );
  INVX0 U902 ( .INP(G7), .ZN(n775) );
  INVX0 U903 ( .INP(n878), .ZN(n870) );
  OA21X1 U904 ( .IN1(n879), .IN2(n880), .IN3(n881), .Q(n861) );
  XOR2X1 U905 ( .IN1(n882), .IN2(keyinput82), .Q(n881) );
  NAND2X0 U906 ( .IN1(n879), .IN2(n880), .QN(n882) );
  XOR2X1 U907 ( .IN1(keyinput63), .IN2(n883), .Q(n880) );
  OA21X1 U908 ( .IN1(G20), .IN2(n884), .IN3(n885), .Q(n883) );
  XOR2X1 U909 ( .IN1(keyinput43), .IN2(n886), .Q(n885) );
  NOR2X0 U910 ( .IN1(G24), .IN2(n887), .QN(n886) );
  INVX0 U911 ( .INP(G24), .ZN(n884) );
  AND2X1 U912 ( .IN1(n888), .IN2(n889), .Q(n879) );
  XOR2X1 U913 ( .IN1(keyinput44), .IN2(n890), .Q(n889) );
  NOR2X0 U914 ( .IN1(n891), .IN2(n578), .QN(n890) );
  XOR2X1 U915 ( .IN1(keyinput45), .IN2(n892), .Q(n888) );
  NOR2X0 U916 ( .IN1(n891), .IN2(n617), .QN(n892) );
  INVX0 U917 ( .INP(G32), .ZN(n617) );
  XOR2X1 U918 ( .IN1(n893), .IN2(keyinput18), .Q(n891) );
  NAND2X0 U919 ( .IN1(G32), .IN2(G28), .QN(n893) );
  INVX0 U920 ( .INP(n649), .ZN(n594) );
  XNOR2X1 U921 ( .IN1(keyinput141), .IN2(n894), .Q(n649) );
  AOI21X1 U922 ( .IN1(n895), .IN2(n896), .IN3(n897), .QN(n894) );
  XNOR2X1 U923 ( .IN1(n898), .IN2(keyinput137), .Q(n897) );
  NAND2X0 U924 ( .IN1(n896), .IN2(n899), .QN(n898) );
  XNOR2X1 U925 ( .IN1(n900), .IN2(keyinput130), .Q(n896) );
  NAND2X0 U926 ( .IN1(n895), .IN2(n899), .QN(n900) );
  NAND2X0 U927 ( .IN1(n901), .IN2(n902), .QN(n899) );
  XOR2X1 U928 ( .IN1(n903), .IN2(keyinput119), .Q(n902) );
  NAND2X0 U929 ( .IN1(n904), .IN2(n905), .QN(n903) );
  XOR2X1 U930 ( .IN1(n906), .IN2(keyinput120), .Q(n901) );
  NAND2X0 U931 ( .IN1(n905), .IN2(n907), .QN(n906) );
  XNOR2X1 U932 ( .IN1(n908), .IN2(keyinput113), .Q(n905) );
  NAND2X0 U933 ( .IN1(n904), .IN2(n907), .QN(n908) );
  XOR2X1 U934 ( .IN1(keyinput107), .IN2(n909), .Q(n907) );
  OA21X1 U935 ( .IN1(n846), .IN2(n910), .IN3(n911), .Q(n909) );
  XOR2X1 U936 ( .IN1(keyinput100), .IN2(n912), .Q(n911) );
  NOR2X0 U937 ( .IN1(n878), .IN2(n910), .QN(n912) );
  XNOR2X1 U938 ( .IN1(n913), .IN2(keyinput96), .Q(n910) );
  OR2X1 U939 ( .IN1(n846), .IN2(n878), .Q(n913) );
  XOR2X1 U940 ( .IN1(n914), .IN2(keyinput86), .Q(n878) );
  NAND2X0 U941 ( .IN1(n915), .IN2(n916), .QN(n914) );
  XOR2X1 U942 ( .IN1(keyinput72), .IN2(n917), .Q(n916) );
  NOR2X0 U943 ( .IN1(n918), .IN2(n919), .QN(n917) );
  XNOR2X1 U944 ( .IN1(keyinput50), .IN2(n920), .Q(n919) );
  XOR2X1 U945 ( .IN1(keyinput73), .IN2(n921), .Q(n915) );
  NOR2X0 U946 ( .IN1(n918), .IN2(n922), .QN(n921) );
  XNOR2X1 U947 ( .IN1(keyinput51), .IN2(n923), .Q(n922) );
  XOR2X1 U948 ( .IN1(n924), .IN2(keyinput64), .Q(n918) );
  NAND2X0 U949 ( .IN1(n925), .IN2(n926), .QN(n924) );
  XOR2X1 U950 ( .IN1(n923), .IN2(keyinput51), .Q(n926) );
  NAND2X0 U951 ( .IN1(n927), .IN2(n928), .QN(n923) );
  XOR2X1 U952 ( .IN1(keyinput25), .IN2(n929), .Q(n928) );
  NOR2X0 U953 ( .IN1(G16), .IN2(n930), .QN(n929) );
  XOR2X1 U954 ( .IN1(n931), .IN2(keyinput26), .Q(n927) );
  NAND2X0 U955 ( .IN1(G16), .IN2(n930), .QN(n931) );
  XOR2X1 U956 ( .IN1(n920), .IN2(keyinput50), .Q(n925) );
  NAND2X0 U957 ( .IN1(n932), .IN2(n933), .QN(n920) );
  XOR2X1 U958 ( .IN1(keyinput23), .IN2(n934), .Q(n933) );
  AND2X1 U959 ( .IN1(n935), .IN2(G13), .Q(n934) );
  XOR2X1 U960 ( .IN1(n936), .IN2(keyinput24), .Q(n932) );
  NAND2X0 U961 ( .IN1(G14), .IN2(n935), .QN(n936) );
  XNOR2X1 U962 ( .IN1(n937), .IN2(keyinput5), .Q(n935) );
  NAND2X0 U963 ( .IN1(G14), .IN2(G13), .QN(n937) );
  XOR2X1 U964 ( .IN1(keyinput85), .IN2(n938), .Q(n846) );
  OA21X1 U965 ( .IN1(n939), .IN2(n940), .IN3(n941), .Q(n938) );
  XOR2X1 U966 ( .IN1(n942), .IN2(keyinput71), .Q(n941) );
  NAND2X0 U967 ( .IN1(n939), .IN2(n940), .QN(n942) );
  XOR3X1 U968 ( .IN1(keyinput49), .IN2(n666), .IN3(n669), .Q(n940) );
  XNOR2X1 U969 ( .IN1(keyinput48), .IN2(n943), .Q(n939) );
  OA21X1 U970 ( .IN1(n944), .IN2(n945), .IN3(n946), .Q(n943) );
  XOR2X1 U971 ( .IN1(keyinput22), .IN2(n947), .Q(n946) );
  NOR2X0 U972 ( .IN1(n758), .IN2(n945), .QN(n947) );
  XNOR2X1 U973 ( .IN1(n948), .IN2(keyinput4), .Q(n945) );
  NAND2X0 U974 ( .IN1(G9), .IN2(G10), .QN(n948) );
  INVX0 U975 ( .INP(G9), .ZN(n944) );
  AND2X1 U976 ( .IN1(G38), .IN2(G41), .Q(n904) );
  XNOR2X1 U977 ( .IN1(n949), .IN2(keyinput93), .Q(n895) );
  NAND2X0 U978 ( .IN1(n950), .IN2(n951), .QN(n949) );
  XOR2X1 U979 ( .IN1(keyinput79), .IN2(n952), .Q(n951) );
  NOR2X0 U980 ( .IN1(n953), .IN2(n954), .QN(n952) );
  XOR2X1 U981 ( .IN1(n955), .IN2(keyinput80), .Q(n950) );
  NAND2X0 U982 ( .IN1(n953), .IN2(n954), .QN(n955) );
  XNOR2X1 U983 ( .IN1(keyinput62), .IN2(n956), .Q(n954) );
  OA21X1 U984 ( .IN1(G30), .IN2(n646), .IN3(n957), .Q(n956) );
  XOR2X1 U985 ( .IN1(n958), .IN2(keyinput41), .Q(n957) );
  NAND2X0 U986 ( .IN1(G30), .IN2(n646), .QN(n958) );
  AOI21X1 U987 ( .IN1(n959), .IN2(G22), .IN3(n960), .QN(n953) );
  XOR2X1 U988 ( .IN1(keyinput40), .IN2(n961), .Q(n960) );
  AND2X1 U989 ( .IN1(G18), .IN2(n959), .Q(n961) );
  XOR2X1 U990 ( .IN1(n962), .IN2(keyinput15), .Q(n959) );
  NAND2X0 U991 ( .IN1(G22), .IN2(G18), .QN(n962) );
  XOR2X1 U992 ( .IN1(n963), .IN2(keyinput164), .Q(n772) );
  NAND3X0 U993 ( .IN1(n964), .IN2(n965), .IN3(n966), .QN(n963) );
  MUX21X1 U994 ( .IN1(n967), .IN2(n968), .S(n696), .Q(n966) );
  NAND3X0 U995 ( .IN1(n969), .IN2(n612), .IN3(n970), .QN(n968) );
  XOR2X1 U996 ( .IN1(n615), .IN2(keyinput143), .Q(n970) );
  XOR2X1 U997 ( .IN1(n703), .IN2(keyinput144), .Q(n969) );
  NAND3X0 U998 ( .IN1(n703), .IN2(n971), .IN3(n972), .QN(n967) );
  XOR2X1 U999 ( .IN1(keyinput145), .IN2(n643), .Q(n972) );
  XOR2X1 U1000 ( .IN1(keyinput146), .IN2(n693), .Q(n971) );
  XNOR2X1 U1001 ( .IN1(n973), .IN2(keyinput158), .Q(n965) );
  NAND3X0 U1002 ( .IN1(n693), .IN2(n696), .IN3(n643), .QN(n973) );
  INVX0 U1003 ( .INP(n615), .ZN(n643) );
  INVX0 U1004 ( .INP(n642), .ZN(n696) );
  XOR2X1 U1005 ( .IN1(n974), .IN2(keyinput159), .Q(n964) );
  NAND4X0 U1006 ( .IN1(n975), .IN2(n976), .IN3(n693), .IN4(n615), .QN(n974) );
  AO22X1 U1007 ( .IN1(n977), .IN2(n978), .IN3(n979), .IN4(n980), .Q(n615) );
  INVX0 U1008 ( .INP(keyinput131), .ZN(n980) );
  NAND2X0 U1009 ( .IN1(n977), .IN2(n981), .QN(n979) );
  AO21X1 U1010 ( .IN1(keyinput131), .IN2(n981), .IN3(n982), .Q(n978) );
  XOR2X1 U1011 ( .IN1(n983), .IN2(keyinput127), .Q(n977) );
  NAND2X0 U1012 ( .IN1(n982), .IN2(n981), .QN(n983) );
  AO22X1 U1013 ( .IN1(n984), .IN2(n985), .IN3(n986), .IN4(n987), .Q(n981) );
  INVX0 U1014 ( .INP(keyinput78), .ZN(n987) );
  NAND2X0 U1015 ( .IN1(n984), .IN2(n988), .QN(n986) );
  AO21X1 U1016 ( .IN1(keyinput78), .IN2(n988), .IN3(n989), .Q(n985) );
  XOR2X1 U1017 ( .IN1(n990), .IN2(keyinput66), .Q(n984) );
  NAND2X0 U1018 ( .IN1(n988), .IN2(n989), .QN(n990) );
  XOR2X1 U1019 ( .IN1(keyinput56), .IN2(n991), .Q(n989) );
  AND2X1 U1020 ( .IN1(n992), .IN2(n993), .Q(n991) );
  XOR2X1 U1021 ( .IN1(keyinput30), .IN2(n994), .Q(n993) );
  NOR2X0 U1022 ( .IN1(G5), .IN2(n995), .QN(n994) );
  XOR2X1 U1023 ( .IN1(n996), .IN2(keyinput31), .Q(n992) );
  NAND2X0 U1024 ( .IN1(G5), .IN2(n995), .QN(n996) );
  INVX0 U1025 ( .INP(G1), .ZN(n995) );
  XNOR2X1 U1026 ( .IN1(keyinput57), .IN2(n997), .Q(n988) );
  OA21X1 U1027 ( .IN1(G9), .IN2(G13), .IN3(n998), .Q(n997) );
  XOR2X1 U1028 ( .IN1(n999), .IN2(keyinput12), .Q(n998) );
  NAND2X0 U1029 ( .IN1(G9), .IN2(G13), .QN(n999) );
  XOR2X1 U1030 ( .IN1(n1000), .IN2(keyinput123), .Q(n982) );
  NAND2X0 U1031 ( .IN1(n1001), .IN2(n1002), .QN(n1000) );
  XOR2X1 U1032 ( .IN1(keyinput116), .IN2(n1003), .Q(n1002) );
  NOR2X0 U1033 ( .IN1(n1004), .IN2(n1005), .QN(n1003) );
  XNOR2X1 U1034 ( .IN1(keyinput110), .IN2(n1006), .Q(n1005) );
  INVX0 U1035 ( .INP(n1007), .ZN(n1004) );
  XOR2X1 U1036 ( .IN1(n1008), .IN2(keyinput115), .Q(n1001) );
  NAND2X0 U1037 ( .IN1(n1009), .IN2(n1007), .QN(n1008) );
  NAND2X0 U1038 ( .IN1(n1009), .IN2(n1010), .QN(n1007) );
  XOR2X1 U1039 ( .IN1(keyinput110), .IN2(n1006), .Q(n1010) );
  AND2X1 U1040 ( .IN1(n1011), .IN2(n1012), .Q(n1006) );
  XOR2X1 U1041 ( .IN1(keyinput103), .IN2(n1013), .Q(n1012) );
  NOR2X0 U1042 ( .IN1(n1014), .IN2(n1015), .QN(n1013) );
  XOR2X1 U1043 ( .IN1(n1016), .IN2(keyinput102), .Q(n1011) );
  NAND2X0 U1044 ( .IN1(n1015), .IN2(n1014), .QN(n1016) );
  AND2X1 U1045 ( .IN1(G33), .IN2(G41), .Q(n1009) );
  INVX0 U1046 ( .INP(n612), .ZN(n693) );
  XNOR2X1 U1047 ( .IN1(keyinput140), .IN2(n1017), .Q(n612) );
  OA21X1 U1048 ( .IN1(n1018), .IN2(n1019), .IN3(n1020), .Q(n1017) );
  XOR2X1 U1049 ( .IN1(n1021), .IN2(keyinput135), .Q(n1020) );
  NAND2X0 U1050 ( .IN1(n1018), .IN2(n1019), .QN(n1021) );
  XNOR3X1 U1051 ( .IN1(keyinput60), .IN2(keyinput59), .IN3(n1022), .Q(n1019)
         );
  XOR2X1 U1052 ( .IN1(n1023), .IN2(n1024), .Q(n1022) );
  OA21X1 U1053 ( .IN1(G4), .IN2(n605), .IN3(n1025), .Q(n1024) );
  XOR2X1 U1054 ( .IN1(n1026), .IN2(keyinput34), .Q(n1025) );
  NAND2X0 U1055 ( .IN1(G4), .IN2(n605), .QN(n1026) );
  INVX0 U1056 ( .INP(G8), .ZN(n605) );
  NAND2X0 U1057 ( .IN1(n1027), .IN2(n1028), .QN(n1023) );
  XOR2X1 U1058 ( .IN1(keyinput35), .IN2(n1029), .Q(n1028) );
  NOR2X0 U1059 ( .IN1(G16), .IN2(n666), .QN(n1029) );
  XOR2X1 U1060 ( .IN1(n1030), .IN2(keyinput36), .Q(n1027) );
  NAND2X0 U1061 ( .IN1(G16), .IN2(n666), .QN(n1030) );
  INVX0 U1062 ( .INP(G12), .ZN(n666) );
  XNOR2X1 U1063 ( .IN1(keyinput125), .IN2(n1031), .Q(n1018) );
  AOI21X1 U1064 ( .IN1(n1032), .IN2(n1033), .IN3(n1034), .QN(n1031) );
  XNOR2X1 U1065 ( .IN1(keyinput117), .IN2(n1035), .Q(n1034) );
  OA21X1 U1066 ( .IN1(n1036), .IN2(n1037), .IN3(n1032), .Q(n1035) );
  XOR2X1 U1067 ( .IN1(keyinput112), .IN2(n1038), .Q(n1032) );
  OA21X1 U1068 ( .IN1(n1036), .IN2(n1037), .IN3(n1033), .Q(n1038) );
  XNOR2X1 U1069 ( .IN1(n1039), .IN2(keyinput1), .Q(n1033) );
  NAND2X0 U1070 ( .IN1(G36), .IN2(G41), .QN(n1039) );
  XNOR2X1 U1071 ( .IN1(n1040), .IN2(keyinput106), .Q(n1037) );
  OR2X1 U1072 ( .IN1(n1041), .IN2(n1015), .Q(n1040) );
  NOR2X0 U1073 ( .IN1(n1042), .IN2(n1041), .QN(n1036) );
  XNOR2X1 U1074 ( .IN1(n1043), .IN2(keyinput98), .Q(n1041) );
  OR2X1 U1075 ( .IN1(n1015), .IN2(n1042), .Q(n1043) );
  XOR2X1 U1076 ( .IN1(n1044), .IN2(keyinput88), .Q(n1015) );
  NAND2X0 U1077 ( .IN1(n1045), .IN2(n1046), .QN(n1044) );
  XOR2X1 U1078 ( .IN1(keyinput75), .IN2(n1047), .Q(n1046) );
  NOR2X0 U1079 ( .IN1(n1048), .IN2(n1049), .QN(n1047) );
  XOR2X1 U1080 ( .IN1(n1050), .IN2(keyinput74), .Q(n1045) );
  NAND2X0 U1081 ( .IN1(n1048), .IN2(n1049), .QN(n1050) );
  XOR2X1 U1082 ( .IN1(keyinput54), .IN2(n1051), .Q(n1049) );
  OA21X1 U1083 ( .IN1(n1052), .IN2(n814), .IN3(n1053), .Q(n1051) );
  XOR2X1 U1084 ( .IN1(keyinput28), .IN2(n1054), .Q(n1053) );
  NOR2X0 U1085 ( .IN1(n1052), .IN2(n595), .QN(n1054) );
  INVX0 U1086 ( .INP(G22), .ZN(n595) );
  INVX0 U1087 ( .INP(G21), .ZN(n814) );
  XOR2X1 U1088 ( .IN1(n1055), .IN2(keyinput8), .Q(n1052) );
  NAND2X0 U1089 ( .IN1(G22), .IN2(G21), .QN(n1055) );
  XOR2X1 U1090 ( .IN1(n836), .IN2(G24), .Q(n1048) );
  INVX0 U1091 ( .INP(G23), .ZN(n836) );
  XOR2X1 U1092 ( .IN1(n642), .IN2(keyinput147), .Q(n976) );
  XNOR2X1 U1093 ( .IN1(keyinput138), .IN2(n1056), .Q(n642) );
  AOI21X1 U1094 ( .IN1(n1057), .IN2(n1058), .IN3(n1059), .QN(n1056) );
  XNOR2X1 U1095 ( .IN1(n1060), .IN2(keyinput132), .Q(n1059) );
  NAND2X0 U1096 ( .IN1(n1058), .IN2(n1061), .QN(n1060) );
  XNOR2X1 U1097 ( .IN1(n1062), .IN2(keyinput128), .Q(n1058) );
  NAND2X0 U1098 ( .IN1(n1061), .IN2(n1057), .QN(n1062) );
  XOR2X1 U1099 ( .IN1(keyinput90), .IN2(n1063), .Q(n1061) );
  OA21X1 U1100 ( .IN1(n1064), .IN2(n1065), .IN3(n1066), .Q(n1063) );
  XOR2X1 U1101 ( .IN1(keyinput67), .IN2(n1067), .Q(n1066) );
  AND2X1 U1102 ( .IN1(n1065), .IN2(n1064), .Q(n1067) );
  XOR2X1 U1103 ( .IN1(G2), .IN2(G6), .Q(n1065) );
  XOR2X1 U1104 ( .IN1(keyinput58), .IN2(n1068), .Q(n1064) );
  OA21X1 U1105 ( .IN1(G14), .IN2(n758), .IN3(n1069), .Q(n1068) );
  XOR2X1 U1106 ( .IN1(n1070), .IN2(keyinput32), .Q(n1069) );
  NAND2X0 U1107 ( .IN1(G14), .IN2(n758), .QN(n1070) );
  INVX0 U1108 ( .INP(G10), .ZN(n758) );
  XNOR3X1 U1109 ( .IN1(keyinput124), .IN2(keyinput111), .IN3(n1071), .Q(n1057)
         );
  XOR2X1 U1110 ( .IN1(n1072), .IN2(n1073), .Q(n1071) );
  NOR2X0 U1111 ( .IN1(n1074), .IN2(n1075), .QN(n1073) );
  XOR2X1 U1112 ( .IN1(keyinput104), .IN2(n1076), .Q(n1075) );
  NOR2X0 U1113 ( .IN1(n1077), .IN2(n1078), .QN(n1076) );
  XOR2X1 U1114 ( .IN1(n1079), .IN2(keyinput105), .Q(n1074) );
  NAND2X0 U1115 ( .IN1(n1077), .IN2(n1078), .QN(n1079) );
  INVX0 U1116 ( .INP(n1042), .ZN(n1078) );
  XNOR2X1 U1117 ( .IN1(keyinput89), .IN2(n1080), .Q(n1042) );
  OA21X1 U1118 ( .IN1(n1081), .IN2(n1082), .IN3(n1083), .Q(n1080) );
  XOR2X1 U1119 ( .IN1(n1084), .IN2(keyinput77), .Q(n1083) );
  NAND2X0 U1120 ( .IN1(n1081), .IN2(n1082), .QN(n1084) );
  AO21X1 U1121 ( .IN1(n635), .IN2(n1085), .IN3(n1086), .Q(n1082) );
  XOR2X1 U1122 ( .IN1(keyinput10), .IN2(n1087), .Q(n1086) );
  NOR2X0 U1123 ( .IN1(n635), .IN2(n1085), .QN(n1087) );
  INVX0 U1124 ( .INP(G30), .ZN(n1085) );
  INVX0 U1125 ( .INP(G29), .ZN(n635) );
  XOR2X1 U1126 ( .IN1(keyinput55), .IN2(n1088), .Q(n1081) );
  OA21X1 U1127 ( .IN1(G32), .IN2(G31), .IN3(n1089), .Q(n1088) );
  XOR2X1 U1128 ( .IN1(n1090), .IN2(keyinput11), .Q(n1089) );
  NAND2X0 U1129 ( .IN1(G31), .IN2(G32), .QN(n1090) );
  INVX0 U1130 ( .INP(n1091), .ZN(n1077) );
  NAND2X0 U1131 ( .IN1(G34), .IN2(G41), .QN(n1072) );
  XOR2X1 U1132 ( .IN1(n703), .IN2(keyinput148), .Q(n975) );
  XOR2X1 U1133 ( .IN1(n1092), .IN2(keyinput139), .Q(n703) );
  NAND2X0 U1134 ( .IN1(n1093), .IN2(n1094), .QN(n1092) );
  XOR2X1 U1135 ( .IN1(keyinput133), .IN2(n1095), .Q(n1094) );
  NOR2X0 U1136 ( .IN1(n1096), .IN2(n1097), .QN(n1095) );
  XOR2X1 U1137 ( .IN1(n1098), .IN2(keyinput134), .Q(n1093) );
  NAND2X0 U1138 ( .IN1(n1096), .IN2(n1097), .QN(n1098) );
  XNOR3X1 U1139 ( .IN1(keyinput0), .IN2(n1099), .IN3(n1100), .Q(n1097) );
  NAND2X0 U1140 ( .IN1(G35), .IN2(G41), .QN(n1100) );
  OA21X1 U1141 ( .IN1(n1014), .IN2(n1091), .IN3(n1101), .Q(n1099) );
  XOR2X1 U1142 ( .IN1(n1102), .IN2(keyinput97), .Q(n1101) );
  NAND2X0 U1143 ( .IN1(n1014), .IN2(n1091), .QN(n1102) );
  NAND2X0 U1144 ( .IN1(n1103), .IN2(n1104), .QN(n1091) );
  NAND3X0 U1145 ( .IN1(n1105), .IN2(n1106), .IN3(n1107), .QN(n1104) );
  XOR2X1 U1146 ( .IN1(keyinput76), .IN2(n1108), .Q(n1103) );
  AND2X1 U1147 ( .IN1(n1105), .IN2(n1109), .Q(n1108) );
  NAND3X0 U1148 ( .IN1(n1106), .IN2(n1109), .IN3(n1107), .QN(n1105) );
  XOR2X1 U1149 ( .IN1(n1110), .IN2(keyinput9), .Q(n1107) );
  NAND2X0 U1150 ( .IN1(G26), .IN2(G25), .QN(n1110) );
  AO21X1 U1151 ( .IN1(G27), .IN2(n578), .IN3(n1111), .Q(n1109) );
  XOR2X1 U1152 ( .IN1(keyinput29), .IN2(n1112), .Q(n1111) );
  NOR2X0 U1153 ( .IN1(G27), .IN2(n578), .QN(n1112) );
  INVX0 U1154 ( .INP(G28), .ZN(n578) );
  NAND2X0 U1155 ( .IN1(n646), .IN2(n651), .QN(n1106) );
  INVX0 U1156 ( .INP(G25), .ZN(n651) );
  INVX0 U1157 ( .INP(G26), .ZN(n646) );
  XNOR2X1 U1158 ( .IN1(keyinput87), .IN2(n1113), .Q(n1014) );
  AOI21X1 U1159 ( .IN1(n1114), .IN2(n1115), .IN3(n1116), .QN(n1113) );
  XNOR2X1 U1160 ( .IN1(keyinput65), .IN2(n1117), .Q(n1116) );
  NOR2X0 U1161 ( .IN1(n1115), .IN2(n1114), .QN(n1117) );
  XOR2X1 U1162 ( .IN1(keyinput52), .IN2(n1118), .Q(n1115) );
  OA21X1 U1163 ( .IN1(G18), .IN2(G17), .IN3(n1119), .Q(n1118) );
  XOR2X1 U1164 ( .IN1(n1120), .IN2(keyinput6), .Q(n1119) );
  NAND2X0 U1165 ( .IN1(G18), .IN2(G17), .QN(n1120) );
  XOR2X1 U1166 ( .IN1(keyinput53), .IN2(n1121), .Q(n1114) );
  OA21X1 U1167 ( .IN1(n707), .IN2(n1122), .IN3(n1123), .Q(n1121) );
  XOR2X1 U1168 ( .IN1(keyinput27), .IN2(n1124), .Q(n1123) );
  NOR2X0 U1169 ( .IN1(n887), .IN2(n1122), .QN(n1124) );
  INVX0 U1170 ( .INP(G20), .ZN(n887) );
  XNOR2X1 U1171 ( .IN1(n1125), .IN2(keyinput7), .Q(n1122) );
  NAND2X0 U1172 ( .IN1(G19), .IN2(G20), .QN(n1125) );
  INVX0 U1173 ( .INP(G19), .ZN(n707) );
  XNOR2X1 U1174 ( .IN1(n1126), .IN2(keyinput91), .Q(n1096) );
  NAND2X0 U1175 ( .IN1(n1127), .IN2(n1128), .QN(n1126) );
  OR3X1 U1176 ( .IN1(n1129), .IN2(n1130), .IN3(n1131), .Q(n1128) );
  XNOR2X1 U1177 ( .IN1(keyinput68), .IN2(n1132), .Q(n1127) );
  OA21X1 U1178 ( .IN1(n1130), .IN2(n1129), .IN3(n1131), .Q(n1132) );
  XOR2X1 U1179 ( .IN1(n669), .IN2(n930), .Q(n1131) );
  INVX0 U1180 ( .INP(G15), .ZN(n930) );
  INVX0 U1181 ( .INP(G11), .ZN(n669) );
  XNOR2X1 U1182 ( .IN1(n1133), .IN2(keyinput33), .Q(n1129) );
  NAND2X0 U1183 ( .IN1(G7), .IN2(n860), .QN(n1133) );
  NOR2X0 U1184 ( .IN1(n860), .IN2(G7), .QN(n1130) );
  INVX0 U1185 ( .INP(G3), .ZN(n860) );
  XOR2X1 U1186 ( .IN1(keyinput236), .IN2(keyinput171), .Q(n790) );
endmodule

