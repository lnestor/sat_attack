
module c880 ( N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, 
        N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, 
        N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, 
        N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, 
        N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, 
        N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, 
        N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73,
         N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106,
         N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152,
         N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207,
         N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268,
         keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5,
         keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11,
         keyinput12, keyinput13, keyinput14, keyinput15, keyinput16,
         keyinput17, keyinput18, keyinput19, keyinput20, keyinput21,
         keyinput22, keyinput23, keyinput24, keyinput25, keyinput26,
         keyinput27, keyinput28, keyinput29, keyinput30, keyinput31,
         keyinput32, keyinput33, keyinput34, keyinput35, keyinput36,
         keyinput37, keyinput38, keyinput39, keyinput40, keyinput41,
         keyinput42, keyinput43, keyinput44, keyinput45, keyinput46,
         keyinput47, keyinput48, keyinput49, keyinput50, keyinput51,
         keyinput52, keyinput53, keyinput54, keyinput55, keyinput56,
         keyinput57, keyinput58, keyinput59, keyinput60, keyinput61,
         keyinput62, keyinput63, keyinput64, keyinput65, keyinput66,
         keyinput67, keyinput68, keyinput69, keyinput70, keyinput71,
         keyinput72, keyinput73, keyinput74, keyinput75, keyinput76,
         keyinput77, keyinput78, keyinput79, keyinput80, keyinput81,
         keyinput82, keyinput83, keyinput84, keyinput85, keyinput86,
         keyinput87, keyinput88, keyinput89, keyinput90, keyinput91,
         keyinput92, keyinput93, keyinput94, keyinput95, keyinput96,
         keyinput97, keyinput98, keyinput99, keyinput100, keyinput101,
         keyinput102, keyinput103, keyinput104, keyinput105, keyinput106,
         keyinput107, keyinput108, keyinput109, keyinput110, keyinput111,
         keyinput112, keyinput113, keyinput114, keyinput115, keyinput116,
         keyinput117, keyinput118, keyinput119, keyinput120, keyinput121,
         keyinput122, keyinput123, keyinput124, keyinput125, keyinput126,
         keyinput127;
  output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446,
         N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866,
         N874, N878, N879, N880;
  wire   n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648;

  XNOR3X1 U346 ( .IN1(keyinput125), .IN2(keyinput124), .IN3(n327), .Q(N878) );
  NAND3X0 U347 ( .IN1(n328), .IN2(n329), .IN3(n330), .QN(n327) );
  OA222X1 U348 ( .IN1(n331), .IN2(n332), .IN3(n333), .IN4(n334), .IN5(n335), 
        .IN6(n336), .Q(n330) );
  XOR2X1 U349 ( .IN1(keyinput121), .IN2(n337), .Q(n329) );
  OA21X1 U350 ( .IN1(n338), .IN2(n339), .IN3(n340), .Q(n337) );
  XOR2X1 U351 ( .IN1(n341), .IN2(keyinput32), .Q(n340) );
  NAND2X0 U352 ( .IN1(N210), .IN2(n342), .QN(n341) );
  XNOR2X1 U353 ( .IN1(keyinput24), .IN2(n343), .Q(n342) );
  XNOR2X1 U354 ( .IN1(keyinput115), .IN2(n344), .Q(n338) );
  OA21X1 U355 ( .IN1(n345), .IN2(n333), .IN3(n346), .Q(n344) );
  XOR2X1 U356 ( .IN1(n347), .IN2(keyinput112), .Q(n346) );
  NAND2X0 U357 ( .IN1(n345), .IN2(n333), .QN(n347) );
  XOR2X1 U358 ( .IN1(n348), .IN2(keyinput74), .Q(n333) );
  NAND2X0 U359 ( .IN1(n349), .IN2(n350), .QN(n348) );
  XOR2X1 U360 ( .IN1(n351), .IN2(keyinput84), .Q(n328) );
  NAND2X0 U361 ( .IN1(N237), .IN2(n352), .QN(n351) );
  XOR2X1 U362 ( .IN1(n353), .IN2(keyinput117), .Q(N865) );
  NAND4X0 U363 ( .IN1(n354), .IN2(n355), .IN3(n356), .IN4(n357), .QN(n353) );
  XOR2X1 U364 ( .IN1(keyinput17), .IN2(n358), .Q(n357) );
  AND2X1 U365 ( .IN1(N116), .IN2(N210), .Q(n358) );
  OA22X1 U366 ( .IN1(n339), .IN2(n359), .IN3(n336), .IN4(n360), .Q(n356) );
  XOR2X1 U367 ( .IN1(keyinput104), .IN2(n361), .Q(n359) );
  MUX21X1 U368 ( .IN1(n362), .IN2(n363), .S(n364), .Q(n361) );
  NAND2X0 U369 ( .IN1(n365), .IN2(n366), .QN(n363) );
  NOR2X0 U370 ( .IN1(n367), .IN2(n368), .QN(n362) );
  XNOR2X1 U371 ( .IN1(n369), .IN2(keyinput81), .Q(n355) );
  AO22X1 U372 ( .IN1(N260), .IN2(N255), .IN3(N246), .IN4(n370), .Q(n369) );
  XNOR2X1 U373 ( .IN1(keyinput100), .IN2(n371), .Q(n354) );
  OA21X1 U374 ( .IN1(n372), .IN2(n373), .IN3(n374), .Q(n371) );
  XOR2X1 U375 ( .IN1(n375), .IN2(keyinput92), .Q(n374) );
  NAND2X0 U376 ( .IN1(n364), .IN2(N228), .QN(n375) );
  AND2X1 U377 ( .IN1(n376), .IN2(n377), .Q(n364) );
  NAND4X0 U378 ( .IN1(n378), .IN2(n379), .IN3(n380), .IN4(n381), .QN(N864) );
  OA222X1 U379 ( .IN1(n336), .IN2(n382), .IN3(n383), .IN4(n372), .IN5(n334), 
        .IN6(n384), .Q(n381) );
  XNOR2X1 U380 ( .IN1(keyinput111), .IN2(n385), .Q(n380) );
  OA22X1 U381 ( .IN1(n386), .IN2(n339), .IN3(n387), .IN4(n388), .Q(n385) );
  INVX0 U382 ( .INP(N111), .ZN(n387) );
  XNOR3X1 U383 ( .IN1(keyinput99), .IN2(n384), .IN3(n389), .Q(n386) );
  NAND3X0 U384 ( .IN1(n390), .IN2(n391), .IN3(n392), .QN(n389) );
  XOR2X1 U385 ( .IN1(keyinput91), .IN2(n373), .Q(n392) );
  XNOR2X1 U386 ( .IN1(keyinput83), .IN2(n393), .Q(n391) );
  XOR2X1 U387 ( .IN1(keyinput94), .IN2(n394), .Q(n390) );
  NAND2X0 U388 ( .IN1(n395), .IN2(n383), .QN(n384) );
  OR2X1 U389 ( .IN1(n396), .IN2(n332), .Q(n379) );
  NAND2X0 U390 ( .IN1(N259), .IN2(N255), .QN(n378) );
  XOR2X1 U391 ( .IN1(n397), .IN2(keyinput120), .Q(N863) );
  NAND3X0 U392 ( .IN1(n398), .IN2(n399), .IN3(n400), .QN(n397) );
  OA222X1 U393 ( .IN1(n401), .IN2(n388), .IN3(n336), .IN4(n402), .IN5(n403), 
        .IN6(n332), .Q(n400) );
  INVX0 U394 ( .INP(N106), .ZN(n401) );
  XOR2X1 U395 ( .IN1(keyinput106), .IN2(n404), .Q(n399) );
  NOR2X0 U396 ( .IN1(n405), .IN2(n339), .QN(n404) );
  XNOR3X1 U397 ( .IN1(keyinput103), .IN2(n406), .IN3(n407), .Q(n405) );
  XNOR2X1 U398 ( .IN1(keyinput98), .IN2(n408), .Q(n398) );
  OA21X1 U399 ( .IN1(n409), .IN2(n372), .IN3(n410), .Q(n408) );
  XOR2X1 U400 ( .IN1(n411), .IN2(keyinput89), .Q(n410) );
  OR2X1 U401 ( .IN1(n334), .IN2(n406), .Q(n411) );
  MUX21X1 U402 ( .IN1(n412), .IN2(n413), .S(keyinput79), .Q(n406) );
  OA21X1 U403 ( .IN1(n403), .IN2(n402), .IN3(n414), .Q(n413) );
  XNOR2X1 U404 ( .IN1(N183), .IN2(n415), .Q(n412) );
  NAND4X0 U405 ( .IN1(n416), .IN2(n417), .IN3(n418), .IN4(n419), .QN(N850) );
  OA22X1 U406 ( .IN1(n339), .IN2(n420), .IN3(n421), .IN4(n334), .Q(n419) );
  INVX0 U407 ( .INP(n422), .ZN(n421) );
  MUX21X1 U408 ( .IN1(n423), .IN2(n424), .S(keyinput93), .Q(n420) );
  XNOR2X1 U409 ( .IN1(n422), .IN2(N261), .Q(n424) );
  NAND2X0 U410 ( .IN1(N261), .IN2(n422), .QN(n423) );
  XNOR2X1 U411 ( .IN1(n425), .IN2(keyinput82), .Q(n422) );
  NAND2X0 U412 ( .IN1(n366), .IN2(n426), .QN(n425) );
  OA22X1 U413 ( .IN1(n336), .IN2(n427), .IN3(n366), .IN4(n372), .Q(n418) );
  INVX0 U414 ( .INP(n367), .ZN(n366) );
  XNOR2X1 U415 ( .IN1(n428), .IN2(keyinput18), .Q(n417) );
  NAND2X0 U416 ( .IN1(N267), .IN2(N255), .QN(n428) );
  OA22X1 U417 ( .IN1(n429), .IN2(n332), .IN3(n430), .IN4(n388), .Q(n416) );
  OA21X1 U418 ( .IN1(n431), .IN2(n432), .IN3(n433), .Q(N768) );
  XOR2X1 U419 ( .IN1(keyinput64), .IN2(n434), .Q(n433) );
  NOR2X0 U420 ( .IN1(n435), .IN2(n436), .QN(n434) );
  XOR2X1 U421 ( .IN1(keyinput62), .IN2(n431), .Q(n436) );
  XOR2X1 U422 ( .IN1(keyinput61), .IN2(n432), .Q(n435) );
  XNOR3X1 U423 ( .IN1(N177), .IN2(N171), .IN3(n437), .Q(n432) );
  XNOR2X1 U424 ( .IN1(N130), .IN2(n438), .Q(n437) );
  OA21X1 U425 ( .IN1(N165), .IN2(N159), .IN3(n439), .Q(n438) );
  XOR2X1 U426 ( .IN1(n440), .IN2(keyinput15), .Q(n439) );
  NAND2X0 U427 ( .IN1(N165), .IN2(N159), .QN(n440) );
  AOI21X1 U428 ( .IN1(n441), .IN2(n442), .IN3(n443), .QN(n431) );
  XOR2X1 U429 ( .IN1(keyinput51), .IN2(n444), .Q(n443) );
  NOR2X0 U430 ( .IN1(n441), .IN2(n442), .QN(n444) );
  INVX0 U431 ( .INP(N207), .ZN(n442) );
  XNOR3X1 U432 ( .IN1(N183), .IN2(n445), .IN3(n446), .Q(n441) );
  XNOR3X1 U433 ( .IN1(keyinput26), .IN2(keyinput25), .IN3(N201), .Q(n446) );
  XNOR2X1 U434 ( .IN1(n360), .IN2(N189), .Q(n445) );
  INVX0 U435 ( .INP(N195), .ZN(n360) );
  OA21X1 U436 ( .IN1(n447), .IN2(n448), .IN3(n449), .Q(N767) );
  XOR2X1 U437 ( .IN1(keyinput63), .IN2(n450), .Q(n449) );
  NOR2X0 U438 ( .IN1(n451), .IN2(n452), .QN(n450) );
  XOR2X1 U439 ( .IN1(keyinput57), .IN2(n447), .Q(n452) );
  INVX0 U440 ( .INP(n448), .ZN(n451) );
  XOR2X1 U441 ( .IN1(keyinput53), .IN2(n453), .Q(n448) );
  OA21X1 U442 ( .IN1(n454), .IN2(n455), .IN3(n456), .Q(n453) );
  XOR2X1 U443 ( .IN1(n457), .IN2(keyinput46), .Q(n456) );
  NAND2X0 U444 ( .IN1(n454), .IN2(n455), .QN(n457) );
  INVX0 U445 ( .INP(N135), .ZN(n455) );
  MUX21X1 U446 ( .IN1(n458), .IN2(n459), .S(n460), .Q(n454) );
  OA21X1 U447 ( .IN1(n461), .IN2(n430), .IN3(n462), .Q(n460) );
  XOR2X1 U448 ( .IN1(n463), .IN2(keyinput12), .Q(n462) );
  NAND2X0 U449 ( .IN1(n461), .IN2(n430), .QN(n463) );
  INVX0 U450 ( .INP(N121), .ZN(n430) );
  INVX0 U451 ( .INP(N126), .ZN(n461) );
  XNOR2X1 U452 ( .IN1(keyinput31), .IN2(n458), .Q(n459) );
  XOR3X1 U453 ( .IN1(keyinput23), .IN2(N116), .IN3(N111), .Q(n458) );
  AND2X1 U454 ( .IN1(n464), .IN2(n465), .Q(n447) );
  XOR2X1 U455 ( .IN1(keyinput45), .IN2(n466), .Q(n465) );
  NOR2X0 U456 ( .IN1(n467), .IN2(N130), .QN(n466) );
  XOR2X1 U457 ( .IN1(n468), .IN2(keyinput44), .Q(n464) );
  NAND2X0 U458 ( .IN1(n467), .IN2(N130), .QN(n468) );
  AOI21X1 U459 ( .IN1(n469), .IN2(n470), .IN3(n471), .QN(n467) );
  XOR2X1 U460 ( .IN1(keyinput30), .IN2(n472), .Q(n471) );
  NOR2X0 U461 ( .IN1(n469), .IN2(n470), .QN(n472) );
  XNOR3X1 U462 ( .IN1(keyinput21), .IN2(n473), .IN3(N91), .Q(n470) );
  XOR2X1 U463 ( .IN1(n474), .IN2(keyinput22), .Q(n469) );
  NAND2X0 U464 ( .IN1(n475), .IN2(n476), .QN(n474) );
  XOR2X1 U465 ( .IN1(n477), .IN2(keyinput10), .Q(n476) );
  NAND2X0 U466 ( .IN1(N101), .IN2(N106), .QN(n477) );
  XOR2X1 U467 ( .IN1(n478), .IN2(keyinput11), .Q(n475) );
  OR2X1 U468 ( .IN1(N106), .IN2(N101), .Q(n478) );
  XOR2X1 U469 ( .IN1(keyinput28), .IN2(n479), .Q(N449) );
  NOR2X0 U470 ( .IN1(n480), .IN2(n481), .QN(n479) );
  XNOR2X1 U471 ( .IN1(n482), .IN2(keyinput5), .Q(n481) );
  NAND3X0 U472 ( .IN1(N68), .IN2(N59), .IN3(N74), .QN(n482) );
  XOR2X1 U473 ( .IN1(n483), .IN2(keyinput27), .Q(N448) );
  NAND2X0 U474 ( .IN1(n484), .IN2(n485), .QN(n483) );
  INVX0 U475 ( .INP(n480), .ZN(n485) );
  XOR2X1 U476 ( .IN1(n486), .IN2(keyinput4), .Q(n484) );
  NAND2X0 U477 ( .IN1(N68), .IN2(N29), .QN(n486) );
  XOR2X1 U478 ( .IN1(n487), .IN2(keyinput127), .Q(N880) );
  NAND3X0 U479 ( .IN1(n488), .IN2(n489), .IN3(n490), .QN(n487) );
  XNOR2X1 U480 ( .IN1(keyinput97), .IN2(n491), .Q(n490) );
  OA21X1 U481 ( .IN1(n372), .IN2(n492), .IN3(n493), .Q(n491) );
  XOR2X1 U482 ( .IN1(keyinput87), .IN2(n494), .Q(n493) );
  NOR2X0 U483 ( .IN1(n495), .IN2(n334), .QN(n494) );
  INVX0 U484 ( .INP(N228), .ZN(n334) );
  XOR2X1 U485 ( .IN1(keyinput122), .IN2(n496), .Q(n489) );
  OA22X1 U486 ( .IN1(n497), .IN2(n339), .IN3(n473), .IN4(n388), .Q(n496) );
  INVX0 U487 ( .INP(N210), .ZN(n388) );
  INVX0 U488 ( .INP(N96), .ZN(n473) );
  INVX0 U489 ( .INP(N219), .ZN(n339) );
  XNOR2X1 U490 ( .IN1(keyinput116), .IN2(n498), .Q(n497) );
  OA21X1 U491 ( .IN1(n495), .IN2(n499), .IN3(n500), .Q(n498) );
  XOR2X1 U492 ( .IN1(n501), .IN2(keyinput113), .Q(n500) );
  NAND2X0 U493 ( .IN1(n499), .IN2(n495), .QN(n501) );
  XNOR2X1 U494 ( .IN1(keyinput109), .IN2(n502), .Q(n499) );
  AND2X1 U495 ( .IN1(n503), .IN2(n504), .Q(n502) );
  XNOR2X1 U496 ( .IN1(keyinput88), .IN2(n505), .Q(n503) );
  XOR2X1 U497 ( .IN1(n506), .IN2(keyinput76), .Q(n495) );
  NAND2X0 U498 ( .IN1(n492), .IN2(n507), .QN(n506) );
  XOR2X1 U499 ( .IN1(keyinput77), .IN2(n508), .Q(n488) );
  OA22X1 U500 ( .IN1(n336), .IN2(n509), .IN3(n510), .IN4(n332), .Q(n508) );
  XOR2X1 U501 ( .IN1(n511), .IN2(keyinput126), .Q(N879) );
  NAND4X0 U502 ( .IN1(n512), .IN2(n513), .IN3(n514), .IN4(n515), .QN(n511) );
  XOR2X1 U503 ( .IN1(n516), .IN2(keyinput16), .Q(n515) );
  NAND2X0 U504 ( .IN1(N210), .IN2(N91), .QN(n516) );
  OA21X1 U505 ( .IN1(n372), .IN2(n517), .IN3(n518), .Q(n514) );
  XOR2X1 U506 ( .IN1(keyinput75), .IN2(n519), .Q(n518) );
  OA22X1 U507 ( .IN1(n336), .IN2(n520), .IN3(n521), .IN4(n332), .Q(n519) );
  INVX0 U508 ( .INP(N246), .ZN(n332) );
  INVX0 U509 ( .INP(N237), .ZN(n372) );
  XOR2X1 U510 ( .IN1(n522), .IN2(keyinput85), .Q(n513) );
  NAND2X0 U511 ( .IN1(n523), .IN2(N228), .QN(n522) );
  XOR2X1 U512 ( .IN1(n524), .IN2(keyinput119), .Q(n512) );
  NAND2X0 U513 ( .IN1(N219), .IN2(n525), .QN(n524) );
  XNOR3X1 U514 ( .IN1(keyinput108), .IN2(n523), .IN3(n526), .Q(n525) );
  NAND3X0 U515 ( .IN1(n527), .IN2(n528), .IN3(n529), .QN(n526) );
  XOR2X1 U516 ( .IN1(n530), .IN2(keyinput107), .Q(n529) );
  NAND2X0 U517 ( .IN1(n531), .IN2(n507), .QN(n530) );
  XOR2X1 U518 ( .IN1(keyinput96), .IN2(n532), .Q(n528) );
  AND2X1 U519 ( .IN1(n507), .IN2(n533), .Q(n532) );
  XNOR2X1 U520 ( .IN1(keyinput86), .IN2(n534), .Q(n527) );
  NOR2X0 U521 ( .IN1(n535), .IN2(n536), .QN(n523) );
  XOR2X1 U522 ( .IN1(keyinput123), .IN2(n537), .Q(N874) );
  NOR2X0 U523 ( .IN1(n538), .IN2(n539), .QN(n537) );
  AO221X1 U524 ( .IN1(N246), .IN2(n540), .IN3(N210), .IN4(N101), .IN5(n541), 
        .Q(n539) );
  XOR2X1 U525 ( .IN1(n542), .IN2(keyinput52), .Q(n541) );
  OR2X1 U526 ( .IN1(n543), .IN2(n336), .Q(n542) );
  XNOR2X1 U527 ( .IN1(n544), .IN2(keyinput33), .Q(n336) );
  NAND4X0 U528 ( .IN1(N73), .IN2(N72), .IN3(n545), .IN4(N68), .QN(n544) );
  NOR2X0 U529 ( .IN1(n546), .IN2(n480), .QN(n545) );
  XNOR2X1 U530 ( .IN1(n547), .IN2(keyinput3), .Q(n480) );
  NAND4X0 U531 ( .IN1(N13), .IN2(N55), .IN3(N1), .IN4(N8), .QN(n547) );
  AO222X1 U532 ( .IN1(n548), .IN2(N228), .IN3(N219), .IN4(n549), .IN5(n533), 
        .IN6(N237), .Q(n538) );
  XOR2X1 U533 ( .IN1(keyinput110), .IN2(n550), .Q(n549) );
  OA21X1 U534 ( .IN1(n533), .IN2(n504), .IN3(n551), .Q(n550) );
  XOR2X1 U535 ( .IN1(keyinput105), .IN2(n552), .Q(n551) );
  NOR2X0 U536 ( .IN1(n548), .IN2(n553), .QN(n552) );
  AND2X1 U537 ( .IN1(n554), .IN2(n505), .Q(n548) );
  INVX0 U538 ( .INP(n533), .ZN(n505) );
  XOR2X1 U539 ( .IN1(n555), .IN2(keyinput9), .Q(N422) );
  NAND2X0 U540 ( .IN1(N36), .IN2(n556), .QN(n555) );
  INVX0 U541 ( .INP(n546), .ZN(n556) );
  NAND2X0 U542 ( .IN1(N42), .IN2(N59), .QN(n546) );
  NAND2X0 U543 ( .IN1(N80), .IN2(n557), .QN(N420) );
  XNOR2X1 U544 ( .IN1(n558), .IN2(keyinput29), .Q(N450) );
  NAND2X0 U545 ( .IN1(N89), .IN2(n559), .QN(n558) );
  NAND2X0 U546 ( .IN1(n560), .IN2(n561), .QN(N446) );
  XOR2X1 U547 ( .IN1(n562), .IN2(keyinput0), .Q(n560) );
  NAND2X0 U548 ( .IN1(n561), .IN2(n563), .QN(N419) );
  XNOR2X1 U549 ( .IN1(keyinput0), .IN2(n562), .Q(n563) );
  AND3X1 U550 ( .IN1(n564), .IN2(N17), .IN3(N13), .Q(n561) );
  XNOR2X1 U551 ( .IN1(n565), .IN2(keyinput20), .Q(N423) );
  NAND2X0 U552 ( .IN1(N90), .IN2(n559), .QN(n565) );
  OR2X1 U553 ( .IN1(N87), .IN2(N88), .Q(n559) );
  XNOR3X1 U554 ( .IN1(keyinput8), .IN2(keyinput19), .IN3(n566), .Q(N421) );
  NAND3X0 U555 ( .IN1(N80), .IN2(N59), .IN3(N36), .QN(n566) );
  AND2X1 U556 ( .IN1(N86), .IN2(N85), .Q(N391) );
  XNOR2X1 U557 ( .IN1(keyinput6), .IN2(n562), .Q(N390) );
  NAND3X0 U558 ( .IN1(N29), .IN2(N42), .IN3(N36), .QN(n562) );
  AND3X1 U559 ( .IN1(N80), .IN2(N29), .IN3(N36), .Q(N389) );
  AND3X1 U560 ( .IN1(N75), .IN2(N42), .IN3(N29), .Q(N388) );
  AND4X1 U561 ( .IN1(N8), .IN2(N17), .IN3(N1), .IN4(N13), .Q(N418) );
  XOR2X1 U562 ( .IN1(keyinput118), .IN2(n567), .Q(N866) );
  NOR2X0 U563 ( .IN1(n352), .IN2(n568), .QN(n567) );
  XOR2X1 U564 ( .IN1(n569), .IN2(keyinput114), .Q(n568) );
  NAND2X0 U565 ( .IN1(n349), .IN2(n570), .QN(n569) );
  INVX0 U566 ( .INP(n345), .ZN(n570) );
  OA21X1 U567 ( .IN1(n571), .IN2(n535), .IN3(n517), .Q(n345) );
  INVX0 U568 ( .INP(n536), .ZN(n517) );
  NOR2X0 U569 ( .IN1(n520), .IN2(n521), .QN(n536) );
  XNOR2X1 U570 ( .IN1(n572), .IN2(keyinput66), .Q(n535) );
  NAND2X0 U571 ( .IN1(n521), .IN2(n520), .QN(n572) );
  INVX0 U572 ( .INP(N165), .ZN(n520) );
  AND3X1 U573 ( .IN1(n573), .IN2(n574), .IN3(n575), .Q(n521) );
  AOI22X1 U574 ( .IN1(N138), .IN2(N51), .IN3(n576), .IN4(N96), .QN(n575) );
  XNOR2X1 U575 ( .IN1(keyinput40), .IN2(n577), .Q(n574) );
  XOR2X1 U576 ( .IN1(n578), .IN2(keyinput39), .Q(n573) );
  NAND2X0 U577 ( .IN1(N146), .IN2(n579), .QN(n578) );
  NOR2X0 U578 ( .IN1(n580), .IN2(n534), .QN(n571) );
  INVX0 U579 ( .INP(n492), .ZN(n534) );
  XNOR2X1 U580 ( .IN1(n581), .IN2(keyinput67), .Q(n492) );
  NAND2X0 U581 ( .IN1(N171), .IN2(n582), .QN(n581) );
  OA21X1 U582 ( .IN1(n533), .IN2(n531), .IN3(n507), .Q(n580) );
  XNOR2X1 U583 ( .IN1(n583), .IN2(keyinput68), .Q(n507) );
  NAND2X0 U584 ( .IN1(n510), .IN2(n509), .QN(n583) );
  INVX0 U585 ( .INP(N171), .ZN(n509) );
  INVX0 U586 ( .INP(n582), .ZN(n510) );
  NAND3X0 U587 ( .IN1(n584), .IN2(n577), .IN3(n585), .QN(n582) );
  XOR2X1 U588 ( .IN1(n586), .IN2(keyinput41), .Q(n585) );
  NAND2X0 U589 ( .IN1(N149), .IN2(n579), .QN(n586) );
  XNOR2X1 U590 ( .IN1(keyinput55), .IN2(n587), .Q(n584) );
  AOI22X1 U591 ( .IN1(n576), .IN2(N101), .IN3(N138), .IN4(N17), .QN(n587) );
  INVX0 U592 ( .INP(n504), .ZN(n531) );
  NAND2X0 U593 ( .IN1(n554), .IN2(n553), .QN(n504) );
  XNOR2X1 U594 ( .IN1(n588), .IN2(keyinput102), .Q(n553) );
  NAND2X0 U595 ( .IN1(n589), .IN2(n409), .QN(n588) );
  XOR2X1 U596 ( .IN1(n590), .IN2(keyinput78), .Q(n409) );
  NAND2X0 U597 ( .IN1(N183), .IN2(n415), .QN(n590) );
  XOR2X1 U598 ( .IN1(n591), .IN2(keyinput101), .Q(n589) );
  NAND2X0 U599 ( .IN1(n407), .IN2(n414), .QN(n591) );
  NAND2X0 U600 ( .IN1(n403), .IN2(n402), .QN(n414) );
  INVX0 U601 ( .INP(N183), .ZN(n402) );
  INVX0 U602 ( .INP(n415), .ZN(n403) );
  AO221X1 U603 ( .IN1(N143), .IN2(n592), .IN3(N111), .IN4(n576), .IN5(n593), 
        .Q(n415) );
  XNOR2X1 U604 ( .IN1(keyinput42), .IN2(n594), .Q(n593) );
  AO221X1 U605 ( .IN1(n595), .IN2(n596), .IN3(n395), .IN4(n597), .IN5(n598), 
        .Q(n407) );
  XNOR2X1 U606 ( .IN1(keyinput90), .IN2(n383), .Q(n598) );
  OR2X1 U607 ( .IN1(n382), .IN2(n396), .Q(n383) );
  NAND3X0 U608 ( .IN1(n599), .IN2(n393), .IN3(n373), .QN(n597) );
  XOR2X1 U609 ( .IN1(n377), .IN2(keyinput80), .Q(n373) );
  XNOR2X1 U610 ( .IN1(n600), .IN2(keyinput71), .Q(n377) );
  NAND2X0 U611 ( .IN1(N195), .IN2(n370), .QN(n600) );
  NAND2X0 U612 ( .IN1(n368), .IN2(n376), .QN(n393) );
  INVX0 U613 ( .INP(n365), .ZN(n368) );
  NAND2X0 U614 ( .IN1(N261), .IN2(n426), .QN(n365) );
  NAND2X0 U615 ( .IN1(n429), .IN2(n427), .QN(n426) );
  NAND2X0 U616 ( .IN1(keyinput95), .IN2(n394), .QN(n599) );
  INVX0 U617 ( .INP(keyinput95), .ZN(n596) );
  NAND2X0 U618 ( .IN1(n394), .IN2(n395), .QN(n595) );
  XNOR2X1 U619 ( .IN1(n601), .IN2(keyinput70), .Q(n395) );
  NAND2X0 U620 ( .IN1(n396), .IN2(n382), .QN(n601) );
  INVX0 U621 ( .INP(N189), .ZN(n382) );
  XNOR2X1 U622 ( .IN1(n602), .IN2(keyinput60), .Q(n396) );
  NAND3X0 U623 ( .IN1(n603), .IN2(n594), .IN3(n604), .QN(n602) );
  XOR2X1 U624 ( .IN1(keyinput48), .IN2(n605), .Q(n604) );
  AND2X1 U625 ( .IN1(n592), .IN2(N146), .Q(n605) );
  NAND2X0 U626 ( .IN1(N116), .IN2(n576), .QN(n603) );
  AND2X1 U627 ( .IN1(n367), .IN2(n376), .Q(n394) );
  XOR2X1 U628 ( .IN1(n606), .IN2(keyinput72), .Q(n376) );
  OR2X1 U629 ( .IN1(n370), .IN2(N195), .Q(n606) );
  NAND3X0 U630 ( .IN1(n607), .IN2(n608), .IN3(n609), .QN(n370) );
  XOR2X1 U631 ( .IN1(n610), .IN2(keyinput49), .Q(n609) );
  NAND2X0 U632 ( .IN1(N149), .IN2(n592), .QN(n610) );
  NAND2X0 U633 ( .IN1(N121), .IN2(n576), .QN(n608) );
  XOR2X1 U634 ( .IN1(n594), .IN2(keyinput43), .Q(n607) );
  NOR2X0 U635 ( .IN1(n427), .IN2(n429), .QN(n367) );
  AND2X1 U636 ( .IN1(n611), .IN2(n594), .Q(n429) );
  NAND3X0 U637 ( .IN1(n612), .IN2(N55), .IN3(n613), .QN(n594) );
  XNOR2X1 U638 ( .IN1(N268), .IN2(keyinput24), .Q(n613) );
  XOR2X1 U639 ( .IN1(keyinput56), .IN2(n614), .Q(n611) );
  OA21X1 U640 ( .IN1(n615), .IN2(n616), .IN3(n617), .Q(n614) );
  XOR2X1 U641 ( .IN1(n618), .IN2(keyinput50), .Q(n617) );
  NAND2X0 U642 ( .IN1(N126), .IN2(n576), .QN(n618) );
  INVX0 U643 ( .INP(n592), .ZN(n615) );
  NAND2X0 U644 ( .IN1(n619), .IN2(N1), .QN(n592) );
  XOR2X1 U645 ( .IN1(n620), .IN2(keyinput35), .Q(n619) );
  NAND2X0 U646 ( .IN1(n621), .IN2(N17), .QN(n620) );
  INVX0 U647 ( .INP(N201), .ZN(n427) );
  XOR2X1 U648 ( .IN1(n622), .IN2(keyinput69), .Q(n554) );
  NAND2X0 U649 ( .IN1(n623), .IN2(n543), .QN(n622) );
  NOR2X0 U650 ( .IN1(n543), .IN2(n623), .QN(n533) );
  INVX0 U651 ( .INP(n540), .ZN(n623) );
  XNOR2X1 U652 ( .IN1(n624), .IN2(keyinput59), .Q(n540) );
  NAND3X0 U653 ( .IN1(n625), .IN2(n626), .IN3(n627), .QN(n624) );
  XOR2X1 U654 ( .IN1(n628), .IN2(keyinput13), .Q(n627) );
  NAND2X0 U655 ( .IN1(N152), .IN2(N138), .QN(n628) );
  NAND2X0 U656 ( .IN1(N106), .IN2(n576), .QN(n626) );
  XNOR2X1 U657 ( .IN1(keyinput47), .IN2(n629), .Q(n625) );
  OA21X1 U658 ( .IN1(n630), .IN2(n616), .IN3(n577), .Q(n629) );
  INVX0 U659 ( .INP(N153), .ZN(n616) );
  INVX0 U660 ( .INP(N177), .ZN(n543) );
  XNOR2X1 U661 ( .IN1(n631), .IN2(keyinput65), .Q(n349) );
  NAND2X0 U662 ( .IN1(n331), .IN2(n335), .QN(n631) );
  XOR2X1 U663 ( .IN1(n350), .IN2(keyinput73), .Q(n352) );
  OR2X1 U664 ( .IN1(n335), .IN2(n331), .Q(n350) );
  XNOR2X1 U665 ( .IN1(n632), .IN2(keyinput58), .Q(n331) );
  NAND3X0 U666 ( .IN1(n633), .IN2(n634), .IN3(n635), .QN(n632) );
  XNOR2X1 U667 ( .IN1(keyinput54), .IN2(n636), .Q(n635) );
  AOI22X1 U668 ( .IN1(N138), .IN2(N8), .IN3(n576), .IN4(N91), .QN(n636) );
  XNOR2X1 U669 ( .IN1(keyinput36), .IN2(n637), .Q(n576) );
  OA21X1 U670 ( .IN1(n638), .IN2(n639), .IN3(n640), .Q(n637) );
  NAND3X0 U671 ( .IN1(N447), .IN2(n641), .IN3(n642), .QN(n640) );
  XOR2X1 U672 ( .IN1(N42), .IN2(N17), .Q(n641) );
  XOR2X1 U673 ( .IN1(keyinput7), .IN2(n643), .Q(n639) );
  AND2X1 U674 ( .IN1(N42), .IN2(n557), .Q(n643) );
  AND2X1 U675 ( .IN1(N75), .IN2(N59), .Q(n557) );
  XOR2X1 U676 ( .IN1(n644), .IN2(keyinput2), .Q(n638) );
  NAND4X0 U677 ( .IN1(N51), .IN2(N1), .IN3(N17), .IN4(N8), .QN(n644) );
  XOR2X1 U678 ( .IN1(keyinput37), .IN2(n645), .Q(n634) );
  AND2X1 U679 ( .IN1(n579), .IN2(N143), .Q(n645) );
  INVX0 U680 ( .INP(n630), .ZN(n579) );
  XNOR2X1 U681 ( .IN1(n646), .IN2(keyinput34), .Q(n630) );
  NAND2X0 U682 ( .IN1(N55), .IN2(n621), .QN(n646) );
  AND2X1 U683 ( .IN1(N447), .IN2(n647), .Q(n621) );
  XOR2X1 U684 ( .IN1(keyinput14), .IN2(n642), .Q(n647) );
  AND2X1 U685 ( .IN1(N59), .IN2(N156), .Q(n642) );
  XNOR2X1 U686 ( .IN1(keyinput38), .IN2(n577), .Q(n633) );
  NAND3X0 U687 ( .IN1(N17), .IN2(n343), .IN3(n612), .QN(n577) );
  AND4X1 U688 ( .IN1(N80), .IN2(N29), .IN3(N447), .IN4(N75), .Q(n612) );
  XOR2X1 U689 ( .IN1(n648), .IN2(keyinput1), .Q(N447) );
  NAND2X0 U690 ( .IN1(N51), .IN2(n564), .QN(n648) );
  AND2X1 U691 ( .IN1(N26), .IN2(N1), .Q(n564) );
  INVX0 U692 ( .INP(N268), .ZN(n343) );
  INVX0 U693 ( .INP(N159), .ZN(n335) );
endmodule

