
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258;

  XNOR2X1 U666 ( .IN1(G32), .IN2(n634), .Q(G1355) );
  NOR2X0 U667 ( .IN1(n635), .IN2(n636), .QN(n634) );
  XNOR2X1 U668 ( .IN1(G31), .IN2(n637), .Q(G1354) );
  NOR2X0 U669 ( .IN1(n638), .IN2(n636), .QN(n637) );
  XNOR2X1 U670 ( .IN1(G30), .IN2(n639), .Q(G1353) );
  NOR2X0 U671 ( .IN1(n640), .IN2(n636), .QN(n639) );
  XNOR2X1 U672 ( .IN1(G29), .IN2(n641), .Q(G1352) );
  NOR2X0 U673 ( .IN1(n642), .IN2(n636), .QN(n641) );
  XOR2X1 U674 ( .IN1(n643), .IN2(keyinput255), .Q(n636) );
  NAND4X0 U675 ( .IN1(n644), .IN2(n645), .IN3(n646), .IN4(n647), .QN(n643) );
  NOR2X0 U676 ( .IN1(n648), .IN2(n649), .QN(n647) );
  XNOR2X1 U677 ( .IN1(n650), .IN2(n651), .Q(G1351) );
  NAND2X0 U678 ( .IN1(n652), .IN2(n653), .QN(n650) );
  XNOR2X1 U679 ( .IN1(n654), .IN2(n655), .Q(G1350) );
  NAND2X0 U680 ( .IN1(n652), .IN2(n656), .QN(n654) );
  XNOR2X1 U681 ( .IN1(n657), .IN2(n658), .Q(G1349) );
  NAND2X0 U682 ( .IN1(n652), .IN2(n659), .QN(n657) );
  XOR2X1 U683 ( .IN1(n660), .IN2(G25), .Q(G1348) );
  NAND2X0 U684 ( .IN1(n652), .IN2(n661), .QN(n660) );
  XOR2X1 U685 ( .IN1(n662), .IN2(keyinput254), .Q(n652) );
  NAND4X0 U686 ( .IN1(n663), .IN2(n644), .IN3(n645), .IN4(n649), .QN(n662) );
  XNOR2X1 U687 ( .IN1(G24), .IN2(n664), .Q(G1347) );
  NOR2X0 U688 ( .IN1(n635), .IN2(n665), .QN(n664) );
  XNOR2X1 U689 ( .IN1(G23), .IN2(n666), .Q(G1346) );
  NOR2X0 U690 ( .IN1(n638), .IN2(n665), .QN(n666) );
  XNOR2X1 U691 ( .IN1(G22), .IN2(n667), .Q(G1345) );
  NOR2X0 U692 ( .IN1(n640), .IN2(n665), .QN(n667) );
  XNOR2X1 U693 ( .IN1(G21), .IN2(n668), .Q(G1344) );
  NOR2X0 U694 ( .IN1(n642), .IN2(n665), .QN(n668) );
  XOR2X1 U695 ( .IN1(n669), .IN2(keyinput253), .Q(n665) );
  NAND4X0 U696 ( .IN1(n670), .IN2(n671), .IN3(n672), .IN4(n645), .QN(n669) );
  XNOR2X1 U697 ( .IN1(G20), .IN2(n673), .Q(G1343) );
  NOR2X0 U698 ( .IN1(n635), .IN2(n674), .QN(n673) );
  XNOR2X1 U699 ( .IN1(G19), .IN2(n675), .Q(G1342) );
  NOR2X0 U700 ( .IN1(n638), .IN2(n674), .QN(n675) );
  XNOR2X1 U701 ( .IN1(G18), .IN2(n676), .Q(G1341) );
  NOR2X0 U702 ( .IN1(n640), .IN2(n674), .QN(n676) );
  XNOR2X1 U703 ( .IN1(G17), .IN2(n677), .Q(G1340) );
  NOR2X0 U704 ( .IN1(n642), .IN2(n674), .QN(n677) );
  XOR2X1 U705 ( .IN1(n678), .IN2(keyinput252), .Q(n674) );
  NAND4X0 U706 ( .IN1(n645), .IN2(n649), .IN3(n648), .IN4(n679), .QN(n678) );
  NOR2X0 U707 ( .IN1(n644), .IN2(n646), .QN(n679) );
  XNOR2X1 U708 ( .IN1(n680), .IN2(keyinput247), .Q(n645) );
  NAND3X0 U709 ( .IN1(n681), .IN2(n682), .IN3(n683), .QN(n680) );
  OA222X1 U710 ( .IN1(n684), .IN2(n685), .IN3(n686), .IN4(n687), .IN5(
        keyinput244), .IN6(n688), .Q(n683) );
  NOR2X0 U711 ( .IN1(n685), .IN2(n656), .QN(n688) );
  NOR2X0 U712 ( .IN1(n659), .IN2(n685), .QN(n686) );
  INVX0 U713 ( .INP(n689), .ZN(n685) );
  AOI22X1 U714 ( .IN1(n687), .IN2(n640), .IN3(n638), .IN4(keyinput244), .QN(
        n684) );
  INVX0 U715 ( .INP(keyinput243), .ZN(n687) );
  XOR2X1 U716 ( .IN1(n690), .IN2(keyinput245), .Q(n682) );
  NAND2X0 U717 ( .IN1(n691), .IN2(n635), .QN(n690) );
  MUX21X1 U718 ( .IN1(n692), .IN2(n693), .S(keyinput242), .Q(n681) );
  AND2X1 U719 ( .IN1(n642), .IN2(n691), .Q(n693) );
  NAND2X0 U720 ( .IN1(n691), .IN2(n642), .QN(n692) );
  XNOR2X1 U721 ( .IN1(G16), .IN2(n694), .Q(G1339) );
  NOR2X0 U722 ( .IN1(n648), .IN2(n695), .QN(n694) );
  XNOR2X1 U723 ( .IN1(G15), .IN2(n696), .Q(G1338) );
  NOR2X0 U724 ( .IN1(n697), .IN2(n695), .QN(n696) );
  XNOR2X1 U725 ( .IN1(G14), .IN2(n698), .Q(G1337) );
  NOR2X0 U726 ( .IN1(n699), .IN2(n695), .QN(n698) );
  MUX21X1 U727 ( .IN1(n700), .IN2(n701), .S(G13), .Q(G1336) );
  NOR2X0 U728 ( .IN1(n646), .IN2(n695), .QN(n701) );
  OR2X1 U729 ( .IN1(n646), .IN2(n695), .Q(n700) );
  XOR2X1 U730 ( .IN1(n702), .IN2(keyinput251), .Q(n695) );
  NAND4X0 U731 ( .IN1(n703), .IN2(n638), .IN3(n704), .IN4(n642), .QN(n702) );
  NOR2X0 U732 ( .IN1(n635), .IN2(n640), .QN(n704) );
  XNOR2X1 U733 ( .IN1(n705), .IN2(n706), .Q(G1335) );
  NAND2X0 U734 ( .IN1(n707), .IN2(n672), .QN(n705) );
  XOR2X1 U735 ( .IN1(n708), .IN2(G11), .Q(G1334) );
  NAND2X0 U736 ( .IN1(n707), .IN2(n649), .QN(n708) );
  XNOR2X1 U737 ( .IN1(n709), .IN2(n710), .Q(G1333) );
  NAND2X0 U738 ( .IN1(n707), .IN2(n644), .QN(n709) );
  XOR2X1 U739 ( .IN1(n711), .IN2(G9), .Q(G1332) );
  NAND2X0 U740 ( .IN1(n707), .IN2(n670), .QN(n711) );
  XOR2X1 U741 ( .IN1(n712), .IN2(keyinput250), .Q(n707) );
  NAND4X0 U742 ( .IN1(n703), .IN2(n689), .IN3(n656), .IN4(n659), .QN(n712) );
  NOR2X0 U743 ( .IN1(n653), .IN2(n661), .QN(n689) );
  XNOR2X1 U744 ( .IN1(G8), .IN2(n713), .Q(G1331) );
  NOR2X0 U745 ( .IN1(n648), .IN2(n714), .QN(n713) );
  XNOR2X1 U746 ( .IN1(G7), .IN2(n715), .Q(G1330) );
  NOR2X0 U747 ( .IN1(n697), .IN2(n714), .QN(n715) );
  XNOR2X1 U748 ( .IN1(G6), .IN2(n716), .Q(G1329) );
  NOR2X0 U749 ( .IN1(n699), .IN2(n714), .QN(n716) );
  MUX21X1 U750 ( .IN1(n717), .IN2(n718), .S(G5), .Q(G1328) );
  NOR2X0 U751 ( .IN1(n646), .IN2(n714), .QN(n718) );
  OR2X1 U752 ( .IN1(n646), .IN2(n714), .Q(n717) );
  XOR2X1 U753 ( .IN1(n719), .IN2(keyinput249), .Q(n714) );
  NAND4X0 U754 ( .IN1(n703), .IN2(n691), .IN3(n661), .IN4(n653), .QN(n719) );
  NOR2X0 U755 ( .IN1(n656), .IN2(n659), .QN(n691) );
  XNOR2X1 U756 ( .IN1(G4), .IN2(n720), .Q(G1327) );
  NOR2X0 U757 ( .IN1(n648), .IN2(n721), .QN(n720) );
  INVX0 U758 ( .INP(n672), .ZN(n648) );
  XNOR2X1 U759 ( .IN1(G3), .IN2(n722), .Q(G1326) );
  NOR2X0 U760 ( .IN1(n697), .IN2(n721), .QN(n722) );
  XNOR2X1 U761 ( .IN1(G2), .IN2(n723), .Q(G1325) );
  NOR2X0 U762 ( .IN1(n699), .IN2(n721), .QN(n723) );
  MUX21X1 U763 ( .IN1(n724), .IN2(n725), .S(n726), .Q(G1324) );
  OR2X1 U764 ( .IN1(n646), .IN2(n721), .Q(n725) );
  NOR2X0 U765 ( .IN1(n646), .IN2(n721), .QN(n724) );
  XOR2X1 U766 ( .IN1(n727), .IN2(keyinput248), .Q(n721) );
  NAND4X0 U767 ( .IN1(n703), .IN2(n640), .IN3(n728), .IN4(n635), .QN(n727) );
  INVX0 U768 ( .INP(n653), .ZN(n635) );
  XNOR2X1 U769 ( .IN1(n729), .IN2(keyinput235), .Q(n653) );
  NAND2X0 U770 ( .IN1(n730), .IN2(n731), .QN(n729) );
  XOR2X1 U771 ( .IN1(keyinput229), .IN2(n732), .Q(n731) );
  NOR2X0 U772 ( .IN1(n733), .IN2(n734), .QN(n732) );
  XNOR2X1 U773 ( .IN1(keyinput205), .IN2(n735), .Q(n734) );
  INVX0 U774 ( .INP(n736), .ZN(n733) );
  XOR2X1 U775 ( .IN1(n737), .IN2(keyinput228), .Q(n730) );
  NAND2X0 U776 ( .IN1(n738), .IN2(n736), .QN(n737) );
  XNOR2X1 U777 ( .IN1(n739), .IN2(keyinput213), .Q(n736) );
  NAND2X0 U778 ( .IN1(n738), .IN2(n740), .QN(n739) );
  XOR2X1 U779 ( .IN1(keyinput205), .IN2(n735), .Q(n740) );
  AND2X1 U780 ( .IN1(n741), .IN2(n742), .Q(n735) );
  XOR2X1 U781 ( .IN1(keyinput196), .IN2(n743), .Q(n742) );
  NOR2X0 U782 ( .IN1(n744), .IN2(n745), .QN(n743) );
  XOR2X1 U783 ( .IN1(keyinput197), .IN2(n746), .Q(n741) );
  NOR2X0 U784 ( .IN1(n745), .IN2(n747), .QN(n746) );
  XOR2X1 U785 ( .IN1(keyinput169), .IN2(n748), .Q(n747) );
  XNOR2X1 U786 ( .IN1(n749), .IN2(keyinput181), .Q(n745) );
  NAND2X0 U787 ( .IN1(n750), .IN2(n751), .QN(n749) );
  INVX0 U788 ( .INP(n744), .ZN(n751) );
  NAND2X0 U789 ( .IN1(G41), .IN2(G40), .QN(n744) );
  XNOR2X1 U790 ( .IN1(keyinput169), .IN2(n748), .Q(n750) );
  AND2X1 U791 ( .IN1(n752), .IN2(n753), .Q(n748) );
  XOR2X1 U792 ( .IN1(n754), .IN2(keyinput156), .Q(n753) );
  NAND2X0 U793 ( .IN1(n755), .IN2(n756), .QN(n754) );
  XOR2X1 U794 ( .IN1(n757), .IN2(keyinput157), .Q(n752) );
  NAND2X0 U795 ( .IN1(n756), .IN2(n758), .QN(n757) );
  XNOR2X1 U796 ( .IN1(n759), .IN2(keyinput145), .Q(n756) );
  NAND2X0 U797 ( .IN1(n755), .IN2(n758), .QN(n759) );
  XOR2X1 U798 ( .IN1(n760), .IN2(keyinput141), .Q(n738) );
  NAND2X0 U799 ( .IN1(n761), .IN2(n762), .QN(n760) );
  XOR2X1 U800 ( .IN1(n763), .IN2(keyinput125), .Q(n762) );
  NAND2X0 U801 ( .IN1(n764), .IN2(n765), .QN(n763) );
  XOR2X1 U802 ( .IN1(n766), .IN2(keyinput124), .Q(n761) );
  NAND2X0 U803 ( .IN1(n764), .IN2(n767), .QN(n766) );
  XOR2X1 U804 ( .IN1(n768), .IN2(keyinput93), .Q(n764) );
  NAND2X0 U805 ( .IN1(n765), .IN2(n767), .QN(n768) );
  XNOR2X1 U806 ( .IN1(n769), .IN2(keyinput76), .Q(n767) );
  NAND2X0 U807 ( .IN1(n770), .IN2(n771), .QN(n769) );
  XOR2X1 U808 ( .IN1(keyinput42), .IN2(n772), .Q(n771) );
  NOR2X0 U809 ( .IN1(G24), .IN2(n773), .QN(n772) );
  XOR2X1 U810 ( .IN1(keyinput43), .IN2(n774), .Q(n770) );
  NOR2X0 U811 ( .IN1(G20), .IN2(n775), .QN(n774) );
  XOR2X1 U812 ( .IN1(n776), .IN2(keyinput77), .Q(n765) );
  NAND2X0 U813 ( .IN1(n777), .IN2(n778), .QN(n776) );
  XOR2X1 U814 ( .IN1(keyinput44), .IN2(n779), .Q(n778) );
  NOR2X0 U815 ( .IN1(G32), .IN2(n651), .QN(n779) );
  XOR2X1 U816 ( .IN1(n780), .IN2(keyinput45), .Q(n777) );
  NAND2X0 U817 ( .IN1(G32), .IN2(n651), .QN(n780) );
  NOR2X0 U818 ( .IN1(n642), .IN2(n638), .QN(n728) );
  INVX0 U819 ( .INP(n656), .ZN(n638) );
  XNOR2X1 U820 ( .IN1(n781), .IN2(keyinput236), .Q(n656) );
  NAND2X0 U821 ( .IN1(n782), .IN2(n783), .QN(n781) );
  XOR2X1 U822 ( .IN1(keyinput227), .IN2(n784), .Q(n783) );
  NOR2X0 U823 ( .IN1(n785), .IN2(n786), .QN(n784) );
  XNOR2X1 U824 ( .IN1(keyinput204), .IN2(n787), .Q(n785) );
  XOR2X1 U825 ( .IN1(n788), .IN2(keyinput226), .Q(n782) );
  NAND2X0 U826 ( .IN1(n789), .IN2(n790), .QN(n788) );
  INVX0 U827 ( .INP(n786), .ZN(n789) );
  XNOR2X1 U828 ( .IN1(n791), .IN2(keyinput212), .Q(n786) );
  NAND2X0 U829 ( .IN1(n792), .IN2(n790), .QN(n791) );
  XNOR2X1 U830 ( .IN1(n793), .IN2(keyinput140), .Q(n790) );
  NAND2X0 U831 ( .IN1(n794), .IN2(n795), .QN(n793) );
  XOR2X1 U832 ( .IN1(keyinput122), .IN2(n796), .Q(n795) );
  NOR2X0 U833 ( .IN1(n797), .IN2(n798), .QN(n796) );
  XNOR2X1 U834 ( .IN1(keyinput74), .IN2(n799), .Q(n798) );
  INVX0 U835 ( .INP(n800), .ZN(n797) );
  XOR2X1 U836 ( .IN1(n801), .IN2(keyinput123), .Q(n794) );
  NAND2X0 U837 ( .IN1(n802), .IN2(n800), .QN(n801) );
  XNOR2X1 U838 ( .IN1(n803), .IN2(keyinput92), .Q(n800) );
  NAND2X0 U839 ( .IN1(n802), .IN2(n804), .QN(n803) );
  XOR2X1 U840 ( .IN1(keyinput74), .IN2(n799), .Q(n804) );
  AND2X1 U841 ( .IN1(n805), .IN2(n806), .Q(n799) );
  XOR2X1 U842 ( .IN1(keyinput38), .IN2(n807), .Q(n806) );
  NOR2X0 U843 ( .IN1(G23), .IN2(n808), .QN(n807) );
  XOR2X1 U844 ( .IN1(keyinput39), .IN2(n809), .Q(n805) );
  AND2X1 U845 ( .IN1(n808), .IN2(G23), .Q(n809) );
  XOR2X1 U846 ( .IN1(n810), .IN2(keyinput75), .Q(n802) );
  NAND2X0 U847 ( .IN1(n811), .IN2(n812), .QN(n810) );
  XOR2X1 U848 ( .IN1(n813), .IN2(keyinput40), .Q(n812) );
  OR2X1 U849 ( .IN1(n655), .IN2(G31), .Q(n813) );
  XOR2X1 U850 ( .IN1(n814), .IN2(keyinput41), .Q(n811) );
  NAND2X0 U851 ( .IN1(G31), .IN2(n655), .QN(n814) );
  XOR2X1 U852 ( .IN1(keyinput204), .IN2(n787), .Q(n792) );
  AND2X1 U853 ( .IN1(n815), .IN2(n816), .Q(n787) );
  XOR2X1 U854 ( .IN1(keyinput194), .IN2(n817), .Q(n816) );
  NOR2X0 U855 ( .IN1(n818), .IN2(n819), .QN(n817) );
  XOR2X1 U856 ( .IN1(keyinput195), .IN2(n820), .Q(n815) );
  NOR2X0 U857 ( .IN1(n818), .IN2(n821), .QN(n820) );
  XOR2X1 U858 ( .IN1(n822), .IN2(keyinput168), .Q(n821) );
  XOR2X1 U859 ( .IN1(n823), .IN2(keyinput180), .Q(n818) );
  NAND2X0 U860 ( .IN1(n824), .IN2(n825), .QN(n823) );
  XNOR2X1 U861 ( .IN1(keyinput168), .IN2(n822), .Q(n825) );
  NAND2X0 U862 ( .IN1(n826), .IN2(n827), .QN(n822) );
  XOR2X1 U863 ( .IN1(n828), .IN2(keyinput154), .Q(n827) );
  NAND2X0 U864 ( .IN1(n829), .IN2(n830), .QN(n828) );
  XOR2X1 U865 ( .IN1(n831), .IN2(keyinput155), .Q(n826) );
  NAND2X0 U866 ( .IN1(n829), .IN2(n832), .QN(n831) );
  XNOR2X1 U867 ( .IN1(n833), .IN2(keyinput144), .Q(n829) );
  NAND2X0 U868 ( .IN1(n832), .IN2(n830), .QN(n833) );
  INVX0 U869 ( .INP(n819), .ZN(n824) );
  NAND2X0 U870 ( .IN1(G39), .IN2(G41), .QN(n819) );
  INVX0 U871 ( .INP(n661), .ZN(n642) );
  XNOR2X1 U872 ( .IN1(n834), .IN2(keyinput237), .Q(n661) );
  NAND2X0 U873 ( .IN1(n835), .IN2(n836), .QN(n834) );
  XOR2X1 U874 ( .IN1(keyinput223), .IN2(n837), .Q(n836) );
  NOR2X0 U875 ( .IN1(n838), .IN2(n839), .QN(n837) );
  XOR2X1 U876 ( .IN1(n840), .IN2(keyinput202), .Q(n839) );
  INVX0 U877 ( .INP(n841), .ZN(n838) );
  XOR2X1 U878 ( .IN1(n842), .IN2(keyinput222), .Q(n835) );
  NAND2X0 U879 ( .IN1(n843), .IN2(n841), .QN(n842) );
  XNOR2X1 U880 ( .IN1(n844), .IN2(keyinput210), .Q(n841) );
  NAND2X0 U881 ( .IN1(n843), .IN2(n845), .QN(n844) );
  XNOR2X1 U882 ( .IN1(keyinput202), .IN2(n840), .Q(n845) );
  NAND2X0 U883 ( .IN1(n846), .IN2(n847), .QN(n840) );
  XNOR2X1 U884 ( .IN1(n848), .IN2(keyinput190), .Q(n847) );
  NAND3X0 U885 ( .IN1(G37), .IN2(G41), .IN3(n849), .QN(n848) );
  XOR2X1 U886 ( .IN1(n850), .IN2(keyinput191), .Q(n846) );
  NAND2X0 U887 ( .IN1(n849), .IN2(n851), .QN(n850) );
  XOR2X1 U888 ( .IN1(n852), .IN2(keyinput178), .Q(n849) );
  NAND3X0 U889 ( .IN1(G41), .IN2(n851), .IN3(G37), .QN(n852) );
  XNOR2X1 U890 ( .IN1(n853), .IN2(keyinput166), .Q(n851) );
  NAND2X0 U891 ( .IN1(n854), .IN2(n855), .QN(n853) );
  XOR2X1 U892 ( .IN1(keyinput150), .IN2(n856), .Q(n855) );
  AND2X1 U893 ( .IN1(n830), .IN2(n857), .Q(n856) );
  XOR2X1 U894 ( .IN1(n858), .IN2(keyinput151), .Q(n854) );
  NAND2X0 U895 ( .IN1(n755), .IN2(n857), .QN(n858) );
  XNOR2X1 U896 ( .IN1(n859), .IN2(keyinput142), .Q(n857) );
  NAND2X0 U897 ( .IN1(n755), .IN2(n830), .QN(n859) );
  XNOR2X1 U898 ( .IN1(n860), .IN2(keyinput126), .Q(n830) );
  NAND2X0 U899 ( .IN1(n861), .IN2(n862), .QN(n860) );
  XOR2X1 U900 ( .IN1(keyinput94), .IN2(n863), .Q(n862) );
  NOR2X0 U901 ( .IN1(n864), .IN2(n865), .QN(n863) );
  XNOR2X1 U902 ( .IN1(keyinput46), .IN2(n866), .Q(n865) );
  XOR2X1 U903 ( .IN1(keyinput95), .IN2(n867), .Q(n861) );
  NOR2X0 U904 ( .IN1(n864), .IN2(n868), .QN(n867) );
  XNOR2X1 U905 ( .IN1(keyinput47), .IN2(n869), .Q(n868) );
  XOR2X1 U906 ( .IN1(n870), .IN2(keyinput78), .Q(n864) );
  NAND2X0 U907 ( .IN1(n871), .IN2(n872), .QN(n870) );
  XOR2X1 U908 ( .IN1(n869), .IN2(keyinput47), .Q(n872) );
  NAND2X0 U909 ( .IN1(n873), .IN2(n874), .QN(n869) );
  XOR2X1 U910 ( .IN1(n875), .IN2(keyinput2), .Q(n874) );
  NAND2X0 U911 ( .IN1(G3), .IN2(n876), .QN(n875) );
  XOR2X1 U912 ( .IN1(n877), .IN2(keyinput3), .Q(n873) );
  OR2X1 U913 ( .IN1(n876), .IN2(G3), .Q(n877) );
  INVX0 U914 ( .INP(G4), .ZN(n876) );
  XOR2X1 U915 ( .IN1(n866), .IN2(keyinput46), .Q(n871) );
  NAND2X0 U916 ( .IN1(n878), .IN2(n879), .QN(n866) );
  XOR2X1 U917 ( .IN1(keyinput0), .IN2(n880), .Q(n879) );
  NOR2X0 U918 ( .IN1(G2), .IN2(n726), .QN(n880) );
  XOR2X1 U919 ( .IN1(n881), .IN2(keyinput1), .Q(n878) );
  NAND2X0 U920 ( .IN1(G2), .IN2(n726), .QN(n881) );
  INVX0 U921 ( .INP(G1), .ZN(n726) );
  XOR2X1 U922 ( .IN1(n882), .IN2(keyinput127), .Q(n755) );
  NAND2X0 U923 ( .IN1(n883), .IN2(n884), .QN(n882) );
  XOR2X1 U924 ( .IN1(n885), .IN2(keyinput97), .Q(n884) );
  NAND2X0 U925 ( .IN1(n886), .IN2(n887), .QN(n885) );
  XOR2X1 U926 ( .IN1(n888), .IN2(keyinput96), .Q(n883) );
  NAND2X0 U927 ( .IN1(n886), .IN2(n889), .QN(n888) );
  XOR2X1 U928 ( .IN1(n890), .IN2(keyinput79), .Q(n886) );
  NAND2X0 U929 ( .IN1(n889), .IN2(n887), .QN(n890) );
  XNOR2X1 U930 ( .IN1(n891), .IN2(keyinput49), .Q(n887) );
  NAND2X0 U931 ( .IN1(n892), .IN2(n893), .QN(n891) );
  XOR2X1 U932 ( .IN1(keyinput6), .IN2(n894), .Q(n893) );
  NOR2X0 U933 ( .IN1(G8), .IN2(n895), .QN(n894) );
  XOR2X1 U934 ( .IN1(keyinput7), .IN2(n896), .Q(n892) );
  AND2X1 U935 ( .IN1(n895), .IN2(G8), .Q(n896) );
  XOR2X1 U936 ( .IN1(n897), .IN2(keyinput48), .Q(n889) );
  NAND2X0 U937 ( .IN1(n898), .IN2(n899), .QN(n897) );
  XOR2X1 U938 ( .IN1(keyinput5), .IN2(n900), .Q(n899) );
  NOR2X0 U939 ( .IN1(G5), .IN2(n901), .QN(n900) );
  XOR2X1 U940 ( .IN1(n902), .IN2(keyinput4), .Q(n898) );
  NAND2X0 U941 ( .IN1(G5), .IN2(n901), .QN(n902) );
  INVX0 U942 ( .INP(G6), .ZN(n901) );
  XOR2X1 U943 ( .IN1(n903), .IN2(keyinput138), .Q(n843) );
  NAND2X0 U944 ( .IN1(n904), .IN2(n905), .QN(n903) );
  XOR2X1 U945 ( .IN1(n906), .IN2(keyinput119), .Q(n905) );
  NAND2X0 U946 ( .IN1(n907), .IN2(n908), .QN(n906) );
  XOR2X1 U947 ( .IN1(n909), .IN2(keyinput118), .Q(n904) );
  NAND2X0 U948 ( .IN1(n907), .IN2(n910), .QN(n909) );
  XOR2X1 U949 ( .IN1(n911), .IN2(keyinput90), .Q(n907) );
  NAND2X0 U950 ( .IN1(n908), .IN2(n910), .QN(n911) );
  XOR3X1 U951 ( .IN1(keyinput70), .IN2(G21), .IN3(G17), .Q(n910) );
  XOR2X1 U952 ( .IN1(n912), .IN2(keyinput71), .Q(n908) );
  NAND2X0 U953 ( .IN1(n913), .IN2(n914), .QN(n912) );
  XOR2X1 U954 ( .IN1(n915), .IN2(keyinput32), .Q(n914) );
  NAND2X0 U955 ( .IN1(G25), .IN2(n916), .QN(n915) );
  XOR2X1 U956 ( .IN1(n917), .IN2(keyinput33), .Q(n913) );
  OR2X1 U957 ( .IN1(n916), .IN2(G25), .Q(n917) );
  INVX0 U958 ( .INP(G29), .ZN(n916) );
  INVX0 U959 ( .INP(n659), .ZN(n640) );
  XNOR2X1 U960 ( .IN1(n918), .IN2(keyinput234), .Q(n659) );
  NAND2X0 U961 ( .IN1(n919), .IN2(n920), .QN(n918) );
  XOR2X1 U962 ( .IN1(keyinput225), .IN2(n921), .Q(n920) );
  NOR2X0 U963 ( .IN1(n922), .IN2(n923), .QN(n921) );
  XOR2X1 U964 ( .IN1(n924), .IN2(keyinput203), .Q(n922) );
  XOR2X1 U965 ( .IN1(n925), .IN2(keyinput224), .Q(n919) );
  NAND2X0 U966 ( .IN1(n926), .IN2(n927), .QN(n925) );
  INVX0 U967 ( .INP(n923), .ZN(n926) );
  XNOR2X1 U968 ( .IN1(n928), .IN2(keyinput211), .Q(n923) );
  NAND2X0 U969 ( .IN1(n929), .IN2(n927), .QN(n928) );
  XNOR2X1 U970 ( .IN1(n930), .IN2(keyinput139), .Q(n927) );
  NAND2X0 U971 ( .IN1(n931), .IN2(n932), .QN(n930) );
  XOR2X1 U972 ( .IN1(keyinput121), .IN2(n933), .Q(n932) );
  NOR2X0 U973 ( .IN1(n934), .IN2(n935), .QN(n933) );
  XOR2X1 U974 ( .IN1(keyinput73), .IN2(n936), .Q(n935) );
  INVX0 U975 ( .INP(n937), .ZN(n934) );
  XOR2X1 U976 ( .IN1(n938), .IN2(keyinput120), .Q(n931) );
  NAND2X0 U977 ( .IN1(n939), .IN2(n937), .QN(n938) );
  XNOR2X1 U978 ( .IN1(n940), .IN2(keyinput91), .Q(n937) );
  NAND2X0 U979 ( .IN1(n941), .IN2(n939), .QN(n940) );
  XNOR2X1 U980 ( .IN1(keyinput73), .IN2(n936), .Q(n941) );
  AND2X1 U981 ( .IN1(n942), .IN2(n943), .Q(n936) );
  XOR2X1 U982 ( .IN1(keyinput36), .IN2(n944), .Q(n943) );
  NOR2X0 U983 ( .IN1(G30), .IN2(n658), .QN(n944) );
  XOR2X1 U984 ( .IN1(keyinput37), .IN2(n945), .Q(n942) );
  NOR2X0 U985 ( .IN1(G26), .IN2(n946), .QN(n945) );
  XOR2X1 U986 ( .IN1(n947), .IN2(keyinput72), .Q(n939) );
  NAND2X0 U987 ( .IN1(n948), .IN2(n949), .QN(n947) );
  XOR2X1 U988 ( .IN1(keyinput34), .IN2(n950), .Q(n949) );
  NOR2X0 U989 ( .IN1(G22), .IN2(n951), .QN(n950) );
  XOR2X1 U990 ( .IN1(keyinput35), .IN2(n952), .Q(n948) );
  NOR2X0 U991 ( .IN1(G18), .IN2(n953), .QN(n952) );
  XNOR2X1 U992 ( .IN1(keyinput203), .IN2(n924), .Q(n929) );
  NAND2X0 U993 ( .IN1(n954), .IN2(n955), .QN(n924) );
  XOR2X1 U994 ( .IN1(keyinput193), .IN2(n956), .Q(n955) );
  NOR2X0 U995 ( .IN1(n957), .IN2(n958), .QN(n956) );
  XOR2X1 U996 ( .IN1(n959), .IN2(keyinput167), .Q(n957) );
  XOR2X1 U997 ( .IN1(n960), .IN2(keyinput192), .Q(n954) );
  NAND2X0 U998 ( .IN1(n961), .IN2(n962), .QN(n960) );
  INVX0 U999 ( .INP(n958), .ZN(n961) );
  XNOR2X1 U1000 ( .IN1(n963), .IN2(keyinput179), .Q(n958) );
  NAND2X0 U1001 ( .IN1(n962), .IN2(n964), .QN(n963) );
  XNOR2X1 U1002 ( .IN1(keyinput167), .IN2(n959), .Q(n964) );
  NAND2X0 U1003 ( .IN1(n965), .IN2(n966), .QN(n959) );
  XOR2X1 U1004 ( .IN1(keyinput152), .IN2(n967), .Q(n966) );
  AND2X1 U1005 ( .IN1(n832), .IN2(n968), .Q(n967) );
  XOR2X1 U1006 ( .IN1(n969), .IN2(keyinput153), .Q(n965) );
  NAND2X0 U1007 ( .IN1(n968), .IN2(n758), .QN(n969) );
  XOR2X1 U1008 ( .IN1(n970), .IN2(keyinput143), .Q(n968) );
  NAND2X0 U1009 ( .IN1(n832), .IN2(n758), .QN(n970) );
  XNOR2X1 U1010 ( .IN1(n971), .IN2(keyinput129), .Q(n758) );
  NAND2X0 U1011 ( .IN1(n972), .IN2(n973), .QN(n971) );
  XOR2X1 U1012 ( .IN1(keyinput100), .IN2(n974), .Q(n973) );
  NOR2X0 U1013 ( .IN1(n975), .IN2(n976), .QN(n974) );
  XOR2X1 U1014 ( .IN1(n977), .IN2(keyinput52), .Q(n975) );
  XOR2X1 U1015 ( .IN1(keyinput101), .IN2(n978), .Q(n972) );
  NOR2X0 U1016 ( .IN1(n979), .IN2(n976), .QN(n978) );
  XNOR2X1 U1017 ( .IN1(n980), .IN2(keyinput81), .Q(n976) );
  NAND2X0 U1018 ( .IN1(n981), .IN2(n982), .QN(n980) );
  XNOR2X1 U1019 ( .IN1(keyinput52), .IN2(n977), .Q(n982) );
  NAND2X0 U1020 ( .IN1(n983), .IN2(n984), .QN(n977) );
  XOR2X1 U1021 ( .IN1(keyinput13), .IN2(n985), .Q(n984) );
  NOR2X0 U1022 ( .IN1(G13), .IN2(n986), .QN(n985) );
  XOR2X1 U1023 ( .IN1(n987), .IN2(keyinput12), .Q(n983) );
  NAND2X0 U1024 ( .IN1(G13), .IN2(n986), .QN(n987) );
  INVX0 U1025 ( .INP(G14), .ZN(n986) );
  XNOR2X1 U1026 ( .IN1(keyinput53), .IN2(n988), .Q(n981) );
  XOR2X1 U1027 ( .IN1(n988), .IN2(keyinput53), .Q(n979) );
  NAND2X0 U1028 ( .IN1(n989), .IN2(n990), .QN(n988) );
  XOR2X1 U1029 ( .IN1(keyinput14), .IN2(n991), .Q(n990) );
  NOR2X0 U1030 ( .IN1(G16), .IN2(n992), .QN(n991) );
  XOR2X1 U1031 ( .IN1(n993), .IN2(keyinput15), .Q(n989) );
  NAND2X0 U1032 ( .IN1(G16), .IN2(n992), .QN(n993) );
  INVX0 U1033 ( .INP(G15), .ZN(n992) );
  XNOR2X1 U1034 ( .IN1(n994), .IN2(keyinput128), .Q(n832) );
  NAND2X0 U1035 ( .IN1(n995), .IN2(n996), .QN(n994) );
  XOR2X1 U1036 ( .IN1(n997), .IN2(keyinput99), .Q(n996) );
  NAND2X0 U1037 ( .IN1(n998), .IN2(n999), .QN(n997) );
  XOR2X1 U1038 ( .IN1(n1000), .IN2(keyinput98), .Q(n995) );
  NAND2X0 U1039 ( .IN1(n998), .IN2(n1001), .QN(n1000) );
  XNOR2X1 U1040 ( .IN1(n1002), .IN2(keyinput80), .Q(n998) );
  NAND2X0 U1041 ( .IN1(n1001), .IN2(n999), .QN(n1002) );
  XNOR2X1 U1042 ( .IN1(n1003), .IN2(keyinput51), .Q(n999) );
  NAND2X0 U1043 ( .IN1(n1004), .IN2(n1005), .QN(n1003) );
  XOR2X1 U1044 ( .IN1(keyinput11), .IN2(n1006), .Q(n1005) );
  NOR2X0 U1045 ( .IN1(G11), .IN2(n706), .QN(n1006) );
  XOR2X1 U1046 ( .IN1(n1007), .IN2(keyinput10), .Q(n1004) );
  NAND2X0 U1047 ( .IN1(G11), .IN2(n706), .QN(n1007) );
  XNOR2X1 U1048 ( .IN1(n1008), .IN2(keyinput50), .Q(n1001) );
  NAND2X0 U1049 ( .IN1(n1009), .IN2(n1010), .QN(n1008) );
  XOR2X1 U1050 ( .IN1(keyinput8), .IN2(n1011), .Q(n1010) );
  AND2X1 U1051 ( .IN1(n710), .IN2(G9), .Q(n1011) );
  XOR2X1 U1052 ( .IN1(keyinput9), .IN2(n1012), .Q(n1009) );
  NOR2X0 U1053 ( .IN1(G9), .IN2(n710), .QN(n1012) );
  AND2X1 U1054 ( .IN1(G38), .IN2(G41), .Q(n962) );
  XOR2X1 U1055 ( .IN1(n1013), .IN2(keyinput246), .Q(n703) );
  NAND3X0 U1056 ( .IN1(n1014), .IN2(n1015), .IN3(n1016), .QN(n1013) );
  OA222X1 U1057 ( .IN1(n1017), .IN2(n1018), .IN3(n1019), .IN4(n1020), .IN5(
        keyinput240), .IN6(n1021), .Q(n1016) );
  NOR2X0 U1058 ( .IN1(n649), .IN2(n1018), .QN(n1021) );
  NOR2X0 U1059 ( .IN1(n1018), .IN2(n644), .QN(n1019) );
  INVX0 U1060 ( .INP(n663), .ZN(n1018) );
  NOR2X0 U1061 ( .IN1(n672), .IN2(n670), .QN(n663) );
  AOI22X1 U1062 ( .IN1(n1020), .IN2(n699), .IN3(n697), .IN4(keyinput240), .QN(
        n1017) );
  INVX0 U1063 ( .INP(n649), .ZN(n697) );
  INVX0 U1064 ( .INP(n644), .ZN(n699) );
  INVX0 U1065 ( .INP(keyinput239), .ZN(n1020) );
  XOR2X1 U1066 ( .IN1(keyinput241), .IN2(n1022), .Q(n1015) );
  NOR2X0 U1067 ( .IN1(n672), .IN2(n1023), .QN(n1022) );
  XNOR2X1 U1068 ( .IN1(n1024), .IN2(keyinput233), .Q(n672) );
  NAND2X0 U1069 ( .IN1(n1025), .IN2(n1026), .QN(n1024) );
  XOR2X1 U1070 ( .IN1(keyinput221), .IN2(n1027), .Q(n1026) );
  NOR2X0 U1071 ( .IN1(n1028), .IN2(n1029), .QN(n1027) );
  XOR2X1 U1072 ( .IN1(n1030), .IN2(keyinput201), .Q(n1028) );
  XOR2X1 U1073 ( .IN1(n1031), .IN2(keyinput220), .Q(n1025) );
  NAND2X0 U1074 ( .IN1(n1032), .IN2(n1033), .QN(n1031) );
  INVX0 U1075 ( .INP(n1029), .ZN(n1032) );
  XNOR2X1 U1076 ( .IN1(n1034), .IN2(keyinput209), .Q(n1029) );
  NAND2X0 U1077 ( .IN1(n1033), .IN2(n1035), .QN(n1034) );
  XNOR2X1 U1078 ( .IN1(keyinput201), .IN2(n1030), .Q(n1035) );
  NAND2X0 U1079 ( .IN1(n1036), .IN2(n1037), .QN(n1030) );
  XOR2X1 U1080 ( .IN1(n1038), .IN2(keyinput189), .Q(n1037) );
  NAND2X0 U1081 ( .IN1(n1039), .IN2(n1040), .QN(n1038) );
  XOR2X1 U1082 ( .IN1(n1041), .IN2(keyinput188), .Q(n1036) );
  NAND3X0 U1083 ( .IN1(G36), .IN2(G41), .IN3(n1039), .QN(n1041) );
  XOR2X1 U1084 ( .IN1(n1042), .IN2(keyinput177), .Q(n1039) );
  NAND3X0 U1085 ( .IN1(G41), .IN2(n1040), .IN3(G36), .QN(n1042) );
  XNOR2X1 U1086 ( .IN1(n1043), .IN2(keyinput173), .Q(n1040) );
  NAND2X0 U1087 ( .IN1(n1044), .IN2(n1045), .QN(n1043) );
  XOR2X1 U1088 ( .IN1(keyinput164), .IN2(n1046), .Q(n1045) );
  NOR2X0 U1089 ( .IN1(n1047), .IN2(n1048), .QN(n1046) );
  INVX0 U1090 ( .INP(n1049), .ZN(n1047) );
  XOR2X1 U1091 ( .IN1(n1050), .IN2(keyinput165), .Q(n1044) );
  OR2X1 U1092 ( .IN1(n1048), .IN2(n1051), .Q(n1050) );
  XNOR2X1 U1093 ( .IN1(n1052), .IN2(keyinput149), .Q(n1048) );
  NAND2X0 U1094 ( .IN1(n1049), .IN2(n1053), .QN(n1052) );
  XOR2X1 U1095 ( .IN1(n1054), .IN2(keyinput137), .Q(n1033) );
  NAND2X0 U1096 ( .IN1(n1055), .IN2(n1056), .QN(n1054) );
  XOR2X1 U1097 ( .IN1(keyinput116), .IN2(n1057), .Q(n1056) );
  NOR2X0 U1098 ( .IN1(n1058), .IN2(n1059), .QN(n1057) );
  XOR2X1 U1099 ( .IN1(keyinput117), .IN2(n1060), .Q(n1055) );
  NOR2X0 U1100 ( .IN1(n1059), .IN2(n1061), .QN(n1060) );
  XOR2X1 U1101 ( .IN1(n1062), .IN2(keyinput89), .Q(n1059) );
  OR2X1 U1102 ( .IN1(n1061), .IN2(n1058), .Q(n1062) );
  XNOR3X1 U1103 ( .IN1(keyinput68), .IN2(G8), .IN3(G4), .Q(n1058) );
  XNOR3X1 U1104 ( .IN1(keyinput69), .IN2(G16), .IN3(n706), .Q(n1061) );
  INVX0 U1105 ( .INP(G12), .ZN(n706) );
  MUX21X1 U1106 ( .IN1(n1063), .IN2(n1064), .S(keyinput238), .Q(n1014) );
  NAND2X0 U1107 ( .IN1(n671), .IN2(n646), .QN(n1064) );
  NOR2X0 U1108 ( .IN1(n670), .IN2(n1023), .QN(n1063) );
  INVX0 U1109 ( .INP(n671), .ZN(n1023) );
  NOR2X0 U1110 ( .IN1(n644), .IN2(n649), .QN(n671) );
  XNOR2X1 U1111 ( .IN1(n1065), .IN2(keyinput232), .Q(n649) );
  NAND2X0 U1112 ( .IN1(n1066), .IN2(n1067), .QN(n1065) );
  XOR2X1 U1113 ( .IN1(keyinput218), .IN2(n1068), .Q(n1067) );
  NOR2X0 U1114 ( .IN1(n1069), .IN2(n1070), .QN(n1068) );
  XOR2X1 U1115 ( .IN1(n1071), .IN2(keyinput136), .Q(n1070) );
  INVX0 U1116 ( .INP(n1072), .ZN(n1069) );
  XOR2X1 U1117 ( .IN1(n1073), .IN2(keyinput219), .Q(n1066) );
  NAND2X0 U1118 ( .IN1(n1074), .IN2(n1072), .QN(n1073) );
  XNOR2X1 U1119 ( .IN1(n1075), .IN2(keyinput208), .Q(n1072) );
  NAND2X0 U1120 ( .IN1(n1074), .IN2(n1076), .QN(n1075) );
  XNOR2X1 U1121 ( .IN1(keyinput136), .IN2(n1071), .Q(n1076) );
  NAND2X0 U1122 ( .IN1(n1077), .IN2(n1078), .QN(n1071) );
  XOR2X1 U1123 ( .IN1(keyinput114), .IN2(n1079), .Q(n1078) );
  AND2X1 U1124 ( .IN1(n1080), .IN2(n1081), .Q(n1079) );
  XOR2X1 U1125 ( .IN1(n1082), .IN2(keyinput115), .Q(n1077) );
  NAND2X0 U1126 ( .IN1(n1081), .IN2(n1083), .QN(n1082) );
  XNOR2X1 U1127 ( .IN1(n1084), .IN2(keyinput88), .Q(n1081) );
  NAND2X0 U1128 ( .IN1(n1083), .IN2(n1080), .QN(n1084) );
  XNOR3X1 U1129 ( .IN1(keyinput66), .IN2(n895), .IN3(G3), .Q(n1080) );
  INVX0 U1130 ( .INP(G7), .ZN(n895) );
  XOR3X1 U1131 ( .IN1(keyinput67), .IN2(G15), .IN3(G11), .Q(n1083) );
  XOR2X1 U1132 ( .IN1(n1085), .IN2(keyinput200), .Q(n1074) );
  NAND2X0 U1133 ( .IN1(n1086), .IN2(n1087), .QN(n1085) );
  XOR2X1 U1134 ( .IN1(keyinput187), .IN2(n1088), .Q(n1087) );
  NOR2X0 U1135 ( .IN1(n1089), .IN2(n1090), .QN(n1088) );
  XNOR2X1 U1136 ( .IN1(keyinput172), .IN2(n1091), .Q(n1090) );
  XOR2X1 U1137 ( .IN1(n1092), .IN2(keyinput186), .Q(n1086) );
  NAND2X0 U1138 ( .IN1(n1093), .IN2(n1094), .QN(n1092) );
  INVX0 U1139 ( .INP(n1089), .ZN(n1093) );
  XNOR2X1 U1140 ( .IN1(n1095), .IN2(keyinput176), .Q(n1089) );
  NAND2X0 U1141 ( .IN1(n1096), .IN2(n1094), .QN(n1095) );
  AND2X1 U1142 ( .IN1(G35), .IN2(G41), .Q(n1094) );
  XOR2X1 U1143 ( .IN1(n1091), .IN2(keyinput172), .Q(n1096) );
  NAND2X0 U1144 ( .IN1(n1097), .IN2(n1098), .QN(n1091) );
  XOR2X1 U1145 ( .IN1(keyinput163), .IN2(n1099), .Q(n1098) );
  AND2X1 U1146 ( .IN1(n1100), .IN2(n1101), .Q(n1099) );
  XOR2X1 U1147 ( .IN1(n1102), .IN2(keyinput162), .Q(n1097) );
  NAND2X0 U1148 ( .IN1(n1100), .IN2(n1103), .QN(n1102) );
  XNOR2X1 U1149 ( .IN1(n1104), .IN2(keyinput148), .Q(n1100) );
  NAND2X0 U1150 ( .IN1(n1101), .IN2(n1103), .QN(n1104) );
  XNOR2X1 U1151 ( .IN1(n1105), .IN2(keyinput231), .Q(n644) );
  NAND2X0 U1152 ( .IN1(n1106), .IN2(n1107), .QN(n1105) );
  XOR2X1 U1153 ( .IN1(keyinput217), .IN2(n1108), .Q(n1107) );
  NOR2X0 U1154 ( .IN1(n1109), .IN2(n1110), .QN(n1108) );
  XNOR2X1 U1155 ( .IN1(keyinput199), .IN2(n1111), .Q(n1109) );
  XOR2X1 U1156 ( .IN1(n1112), .IN2(keyinput216), .Q(n1106) );
  NAND2X0 U1157 ( .IN1(n1113), .IN2(n1114), .QN(n1112) );
  INVX0 U1158 ( .INP(n1110), .ZN(n1113) );
  XNOR2X1 U1159 ( .IN1(n1115), .IN2(keyinput207), .Q(n1110) );
  NAND2X0 U1160 ( .IN1(n1114), .IN2(n1116), .QN(n1115) );
  XOR2X1 U1161 ( .IN1(keyinput199), .IN2(n1111), .Q(n1116) );
  AND2X1 U1162 ( .IN1(n1117), .IN2(n1118), .Q(n1111) );
  XNOR2X1 U1163 ( .IN1(n1119), .IN2(keyinput184), .Q(n1118) );
  NAND3X0 U1164 ( .IN1(G41), .IN2(n1120), .IN3(G34), .QN(n1119) );
  XOR2X1 U1165 ( .IN1(n1121), .IN2(keyinput185), .Q(n1117) );
  NAND2X0 U1166 ( .IN1(n1120), .IN2(n1122), .QN(n1121) );
  XNOR2X1 U1167 ( .IN1(n1123), .IN2(keyinput175), .Q(n1120) );
  NAND3X0 U1168 ( .IN1(G41), .IN2(n1122), .IN3(G34), .QN(n1123) );
  XNOR2X1 U1169 ( .IN1(n1124), .IN2(keyinput171), .Q(n1122) );
  NAND2X0 U1170 ( .IN1(n1125), .IN2(n1126), .QN(n1124) );
  XOR2X1 U1171 ( .IN1(keyinput160), .IN2(n1127), .Q(n1126) );
  NOR2X0 U1172 ( .IN1(n1128), .IN2(n1129), .QN(n1127) );
  XOR2X1 U1173 ( .IN1(keyinput161), .IN2(n1130), .Q(n1125) );
  NOR2X0 U1174 ( .IN1(n1051), .IN2(n1128), .QN(n1130) );
  XOR2X1 U1175 ( .IN1(n1131), .IN2(keyinput147), .Q(n1128) );
  NAND2X0 U1176 ( .IN1(n1101), .IN2(n1053), .QN(n1131) );
  INVX0 U1177 ( .INP(n1129), .ZN(n1101) );
  XNOR2X1 U1178 ( .IN1(n1132), .IN2(keyinput132), .Q(n1129) );
  NAND2X0 U1179 ( .IN1(n1133), .IN2(n1134), .QN(n1132) );
  XOR2X1 U1180 ( .IN1(keyinput106), .IN2(n1135), .Q(n1134) );
  NOR2X0 U1181 ( .IN1(n1136), .IN2(n1137), .QN(n1135) );
  XOR2X1 U1182 ( .IN1(n1138), .IN2(keyinput58), .Q(n1137) );
  XOR2X1 U1183 ( .IN1(keyinput107), .IN2(n1139), .Q(n1133) );
  NOR2X0 U1184 ( .IN1(n1136), .IN2(n1140), .QN(n1139) );
  XNOR2X1 U1185 ( .IN1(keyinput59), .IN2(n1141), .Q(n1140) );
  XOR2X1 U1186 ( .IN1(n1142), .IN2(keyinput84), .Q(n1136) );
  NAND2X0 U1187 ( .IN1(n1143), .IN2(n1144), .QN(n1142) );
  XNOR2X1 U1188 ( .IN1(keyinput58), .IN2(n1138), .Q(n1144) );
  NAND2X0 U1189 ( .IN1(n1145), .IN2(n1146), .QN(n1138) );
  XOR2X1 U1190 ( .IN1(keyinput25), .IN2(n1147), .Q(n1146) );
  NOR2X0 U1191 ( .IN1(G25), .IN2(n658), .QN(n1147) );
  XOR2X1 U1192 ( .IN1(n1148), .IN2(keyinput24), .Q(n1145) );
  NAND2X0 U1193 ( .IN1(G25), .IN2(n658), .QN(n1148) );
  INVX0 U1194 ( .INP(G26), .ZN(n658) );
  XOR2X1 U1195 ( .IN1(n1141), .IN2(keyinput59), .Q(n1143) );
  NAND2X0 U1196 ( .IN1(n1149), .IN2(n1150), .QN(n1141) );
  XOR2X1 U1197 ( .IN1(n1151), .IN2(keyinput26), .Q(n1150) );
  NAND2X0 U1198 ( .IN1(G27), .IN2(n651), .QN(n1151) );
  INVX0 U1199 ( .INP(G28), .ZN(n651) );
  XOR2X1 U1200 ( .IN1(n1152), .IN2(keyinput27), .Q(n1149) );
  NAND2X0 U1201 ( .IN1(G28), .IN2(n655), .QN(n1152) );
  INVX0 U1202 ( .INP(G27), .ZN(n655) );
  INVX0 U1203 ( .INP(n1053), .ZN(n1051) );
  XNOR2X1 U1204 ( .IN1(n1153), .IN2(keyinput133), .Q(n1053) );
  NAND2X0 U1205 ( .IN1(n1154), .IN2(n1155), .QN(n1153) );
  XOR2X1 U1206 ( .IN1(n1156), .IN2(keyinput109), .Q(n1155) );
  NAND2X0 U1207 ( .IN1(n1157), .IN2(n1158), .QN(n1156) );
  XOR2X1 U1208 ( .IN1(n1159), .IN2(keyinput108), .Q(n1154) );
  NAND2X0 U1209 ( .IN1(n1160), .IN2(n1158), .QN(n1159) );
  XNOR2X1 U1210 ( .IN1(n1161), .IN2(keyinput85), .Q(n1158) );
  NAND2X0 U1211 ( .IN1(n1157), .IN2(n1160), .QN(n1161) );
  XOR2X1 U1212 ( .IN1(n1162), .IN2(keyinput61), .Q(n1157) );
  NAND2X0 U1213 ( .IN1(n1163), .IN2(n1164), .QN(n1162) );
  XOR2X1 U1214 ( .IN1(keyinput31), .IN2(n1165), .Q(n1164) );
  NOR2X0 U1215 ( .IN1(G31), .IN2(n1166), .QN(n1165) );
  XOR2X1 U1216 ( .IN1(n1167), .IN2(keyinput30), .Q(n1163) );
  NAND2X0 U1217 ( .IN1(G31), .IN2(n1166), .QN(n1167) );
  INVX0 U1218 ( .INP(G32), .ZN(n1166) );
  XOR2X1 U1219 ( .IN1(n1168), .IN2(keyinput60), .Q(n1160) );
  NAND2X0 U1220 ( .IN1(n1169), .IN2(n1170), .QN(n1168) );
  XOR2X1 U1221 ( .IN1(keyinput29), .IN2(n1171), .Q(n1170) );
  NOR2X0 U1222 ( .IN1(G29), .IN2(n946), .QN(n1171) );
  XOR2X1 U1223 ( .IN1(n1172), .IN2(keyinput28), .Q(n1169) );
  NAND2X0 U1224 ( .IN1(G29), .IN2(n946), .QN(n1172) );
  INVX0 U1225 ( .INP(G30), .ZN(n946) );
  XOR2X1 U1226 ( .IN1(n1173), .IN2(keyinput135), .Q(n1114) );
  NAND2X0 U1227 ( .IN1(n1174), .IN2(n1175), .QN(n1173) );
  XOR2X1 U1228 ( .IN1(keyinput112), .IN2(n1176), .Q(n1175) );
  AND2X1 U1229 ( .IN1(n1177), .IN2(n1178), .Q(n1176) );
  XOR2X1 U1230 ( .IN1(n1179), .IN2(keyinput113), .Q(n1174) );
  NAND2X0 U1231 ( .IN1(n1177), .IN2(n1180), .QN(n1179) );
  XNOR2X1 U1232 ( .IN1(n1181), .IN2(keyinput87), .Q(n1177) );
  NAND2X0 U1233 ( .IN1(n1178), .IN2(n1180), .QN(n1181) );
  XNOR3X1 U1234 ( .IN1(keyinput65), .IN2(G14), .IN3(n710), .Q(n1180) );
  INVX0 U1235 ( .INP(G10), .ZN(n710) );
  XNOR3X1 U1236 ( .IN1(keyinput64), .IN2(G6), .IN3(G2), .Q(n1178) );
  INVX0 U1237 ( .INP(n646), .ZN(n670) );
  XNOR2X1 U1238 ( .IN1(n1182), .IN2(keyinput230), .Q(n646) );
  NAND2X0 U1239 ( .IN1(n1183), .IN2(n1184), .QN(n1182) );
  XOR2X1 U1240 ( .IN1(keyinput214), .IN2(n1185), .Q(n1184) );
  NOR2X0 U1241 ( .IN1(n1186), .IN2(n1187), .QN(n1185) );
  XOR2X1 U1242 ( .IN1(n1188), .IN2(keyinput134), .Q(n1186) );
  XOR2X1 U1243 ( .IN1(keyinput215), .IN2(n1189), .Q(n1183) );
  NOR2X0 U1244 ( .IN1(n1190), .IN2(n1187), .QN(n1189) );
  XNOR2X1 U1245 ( .IN1(n1191), .IN2(keyinput206), .Q(n1187) );
  NAND2X0 U1246 ( .IN1(n1192), .IN2(n1193), .QN(n1191) );
  XNOR2X1 U1247 ( .IN1(keyinput134), .IN2(n1188), .Q(n1193) );
  NAND2X0 U1248 ( .IN1(n1194), .IN2(n1195), .QN(n1188) );
  XOR2X1 U1249 ( .IN1(keyinput110), .IN2(n1196), .Q(n1195) );
  AND2X1 U1250 ( .IN1(n1197), .IN2(n1198), .Q(n1196) );
  XOR2X1 U1251 ( .IN1(n1199), .IN2(keyinput111), .Q(n1194) );
  NAND2X0 U1252 ( .IN1(n1198), .IN2(n1200), .QN(n1199) );
  XOR2X1 U1253 ( .IN1(n1201), .IN2(keyinput86), .Q(n1198) );
  NAND2X0 U1254 ( .IN1(n1197), .IN2(n1200), .QN(n1201) );
  XOR3X1 U1255 ( .IN1(keyinput63), .IN2(G9), .IN3(G13), .Q(n1200) );
  XNOR3X1 U1256 ( .IN1(keyinput62), .IN2(G5), .IN3(G1), .Q(n1197) );
  XNOR2X1 U1257 ( .IN1(keyinput198), .IN2(n1202), .Q(n1192) );
  XOR2X1 U1258 ( .IN1(n1202), .IN2(keyinput198), .Q(n1190) );
  NAND2X0 U1259 ( .IN1(n1203), .IN2(n1204), .QN(n1202) );
  XOR2X1 U1260 ( .IN1(n1205), .IN2(keyinput183), .Q(n1204) );
  NAND2X0 U1261 ( .IN1(n1206), .IN2(n1207), .QN(n1205) );
  XOR2X1 U1262 ( .IN1(n1208), .IN2(keyinput182), .Q(n1203) );
  NAND3X0 U1263 ( .IN1(G41), .IN2(n1206), .IN3(G33), .QN(n1208) );
  XNOR2X1 U1264 ( .IN1(n1209), .IN2(keyinput174), .Q(n1206) );
  NAND3X0 U1265 ( .IN1(G41), .IN2(n1207), .IN3(G33), .QN(n1209) );
  XNOR2X1 U1266 ( .IN1(n1210), .IN2(keyinput170), .Q(n1207) );
  NAND2X0 U1267 ( .IN1(n1211), .IN2(n1212), .QN(n1210) );
  XOR2X1 U1268 ( .IN1(n1213), .IN2(keyinput158), .Q(n1212) );
  NAND2X0 U1269 ( .IN1(n1214), .IN2(n1103), .QN(n1213) );
  XOR2X1 U1270 ( .IN1(n1215), .IN2(keyinput159), .Q(n1211) );
  NAND2X0 U1271 ( .IN1(n1214), .IN2(n1049), .QN(n1215) );
  XOR2X1 U1272 ( .IN1(n1216), .IN2(keyinput146), .Q(n1214) );
  NAND2X0 U1273 ( .IN1(n1049), .IN2(n1103), .QN(n1216) );
  XNOR2X1 U1274 ( .IN1(n1217), .IN2(keyinput130), .Q(n1103) );
  NAND2X0 U1275 ( .IN1(n1218), .IN2(n1219), .QN(n1217) );
  XOR2X1 U1276 ( .IN1(keyinput102), .IN2(n1220), .Q(n1219) );
  NOR2X0 U1277 ( .IN1(n1221), .IN2(n1222), .QN(n1220) );
  XOR2X1 U1278 ( .IN1(n1223), .IN2(keyinput54), .Q(n1221) );
  XOR2X1 U1279 ( .IN1(n1224), .IN2(keyinput103), .Q(n1218) );
  NAND2X0 U1280 ( .IN1(n1225), .IN2(n1226), .QN(n1224) );
  INVX0 U1281 ( .INP(n1222), .ZN(n1225) );
  XNOR2X1 U1282 ( .IN1(n1227), .IN2(keyinput82), .Q(n1222) );
  NAND2X0 U1283 ( .IN1(n1226), .IN2(n1228), .QN(n1227) );
  XNOR2X1 U1284 ( .IN1(keyinput54), .IN2(n1223), .Q(n1228) );
  NAND2X0 U1285 ( .IN1(n1229), .IN2(n1230), .QN(n1223) );
  XOR2X1 U1286 ( .IN1(keyinput17), .IN2(n1231), .Q(n1230) );
  NOR2X0 U1287 ( .IN1(G17), .IN2(n951), .QN(n1231) );
  XOR2X1 U1288 ( .IN1(n1232), .IN2(keyinput16), .Q(n1229) );
  NAND2X0 U1289 ( .IN1(G17), .IN2(n951), .QN(n1232) );
  INVX0 U1290 ( .INP(G18), .ZN(n951) );
  XOR2X1 U1291 ( .IN1(n1233), .IN2(keyinput55), .Q(n1226) );
  NAND2X0 U1292 ( .IN1(n1234), .IN2(n1235), .QN(n1233) );
  XOR2X1 U1293 ( .IN1(keyinput18), .IN2(n1236), .Q(n1235) );
  NOR2X0 U1294 ( .IN1(G20), .IN2(n808), .QN(n1236) );
  INVX0 U1295 ( .INP(G19), .ZN(n808) );
  XOR2X1 U1296 ( .IN1(keyinput19), .IN2(n1237), .Q(n1234) );
  NOR2X0 U1297 ( .IN1(G19), .IN2(n773), .QN(n1237) );
  INVX0 U1298 ( .INP(G20), .ZN(n773) );
  XNOR2X1 U1299 ( .IN1(n1238), .IN2(keyinput131), .Q(n1049) );
  NAND2X0 U1300 ( .IN1(n1239), .IN2(n1240), .QN(n1238) );
  XOR2X1 U1301 ( .IN1(keyinput104), .IN2(n1241), .Q(n1240) );
  NOR2X0 U1302 ( .IN1(n1242), .IN2(n1243), .QN(n1241) );
  XNOR2X1 U1303 ( .IN1(keyinput56), .IN2(n1244), .Q(n1243) );
  INVX0 U1304 ( .INP(n1245), .ZN(n1242) );
  XOR2X1 U1305 ( .IN1(n1246), .IN2(keyinput105), .Q(n1239) );
  NAND2X0 U1306 ( .IN1(n1247), .IN2(n1245), .QN(n1246) );
  XNOR2X1 U1307 ( .IN1(n1248), .IN2(keyinput83), .Q(n1245) );
  NAND2X0 U1308 ( .IN1(n1249), .IN2(n1247), .QN(n1248) );
  XOR2X1 U1309 ( .IN1(n1244), .IN2(keyinput56), .Q(n1249) );
  NAND2X0 U1310 ( .IN1(n1250), .IN2(n1251), .QN(n1244) );
  XOR2X1 U1311 ( .IN1(keyinput21), .IN2(n1252), .Q(n1251) );
  NOR2X0 U1312 ( .IN1(G21), .IN2(n953), .QN(n1252) );
  XOR2X1 U1313 ( .IN1(n1253), .IN2(keyinput20), .Q(n1250) );
  NAND2X0 U1314 ( .IN1(G21), .IN2(n953), .QN(n1253) );
  INVX0 U1315 ( .INP(G22), .ZN(n953) );
  XOR2X1 U1316 ( .IN1(n1254), .IN2(keyinput57), .Q(n1247) );
  NAND2X0 U1317 ( .IN1(n1255), .IN2(n1256), .QN(n1254) );
  XOR2X1 U1318 ( .IN1(keyinput23), .IN2(n1257), .Q(n1256) );
  NOR2X0 U1319 ( .IN1(G23), .IN2(n775), .QN(n1257) );
  XOR2X1 U1320 ( .IN1(n1258), .IN2(keyinput22), .Q(n1255) );
  NAND2X0 U1321 ( .IN1(G23), .IN2(n775), .QN(n1258) );
  INVX0 U1322 ( .INP(G24), .ZN(n775) );
endmodule

