
module c1355 ( G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, 
        G1329, G1330, G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, 
        G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, G1348, 
        G1349, G1350, G1351, G1352, G1353, G1354, G1355, G14, G15, G16, G17, 
        G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
        G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, 
        G7, G8, G9, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21,
         G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34,
         G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333,
         G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343,
         G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353,
         G1354, G1355;
  wire   n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761;

  XOR3X1 U428 ( .IN1(keyinput122), .IN2(keyinput112), .IN3(n401), .Q(G1343) );
  NOR2X0 U429 ( .IN1(n402), .IN2(n403), .QN(n401) );
  XOR2X1 U430 ( .IN1(keyinput99), .IN2(n404), .Q(n403) );
  AND2X1 U431 ( .IN1(n405), .IN2(n406), .Q(n404) );
  XOR2X1 U432 ( .IN1(n407), .IN2(keyinput98), .Q(n402) );
  NAND2X0 U433 ( .IN1(n406), .IN2(G20), .QN(n407) );
  XOR2X1 U434 ( .IN1(n408), .IN2(keyinput89), .Q(n406) );
  NAND2X0 U435 ( .IN1(G20), .IN2(n405), .QN(n408) );
  XNOR2X1 U436 ( .IN1(n409), .IN2(keyinput81), .Q(n405) );
  NAND2X0 U437 ( .IN1(n410), .IN2(n411), .QN(n409) );
  XOR2X1 U438 ( .IN1(n412), .IN2(keyinput120), .Q(G1328) );
  MUX21X1 U439 ( .IN1(n413), .IN2(n414), .S(G5), .Q(n412) );
  NOR2X0 U440 ( .IN1(n415), .IN2(n416), .QN(n414) );
  OR2X1 U441 ( .IN1(n416), .IN2(n415), .Q(n413) );
  MUX21X1 U442 ( .IN1(n417), .IN2(n418), .S(G31), .Q(G1354) );
  NOR2X0 U443 ( .IN1(n419), .IN2(n420), .QN(n418) );
  NAND2X0 U444 ( .IN1(n421), .IN2(n422), .QN(n417) );
  XOR2X1 U445 ( .IN1(n423), .IN2(n424), .Q(G1353) );
  NOR2X0 U446 ( .IN1(n420), .IN2(n425), .QN(n424) );
  XOR2X1 U447 ( .IN1(n426), .IN2(G28), .Q(G1351) );
  NAND2X0 U448 ( .IN1(n427), .IN2(n411), .QN(n426) );
  XOR2X1 U449 ( .IN1(n428), .IN2(G27), .Q(G1350) );
  NAND2X0 U450 ( .IN1(n427), .IN2(n421), .QN(n428) );
  XOR2X1 U451 ( .IN1(n429), .IN2(G26), .Q(G1349) );
  NAND2X0 U452 ( .IN1(n427), .IN2(n430), .QN(n429) );
  XOR2X1 U453 ( .IN1(n431), .IN2(G25), .Q(G1348) );
  NAND2X0 U454 ( .IN1(n427), .IN2(n432), .QN(n431) );
  AND3X1 U455 ( .IN1(n433), .IN2(n415), .IN3(n434), .Q(n427) );
  XOR2X1 U456 ( .IN1(n435), .IN2(G19), .Q(G1342) );
  NAND2X0 U457 ( .IN1(n410), .IN2(n421), .QN(n435) );
  XOR2X1 U458 ( .IN1(n436), .IN2(G18), .Q(G1341) );
  NAND2X0 U459 ( .IN1(n410), .IN2(n430), .QN(n436) );
  XOR2X1 U460 ( .IN1(n437), .IN2(G16), .Q(G1339) );
  NAND2X0 U461 ( .IN1(n438), .IN2(n439), .QN(n437) );
  XOR2X1 U462 ( .IN1(n440), .IN2(G15), .Q(G1338) );
  NAND2X0 U463 ( .IN1(n438), .IN2(n441), .QN(n440) );
  XOR2X1 U464 ( .IN1(n442), .IN2(G14), .Q(G1337) );
  NAND2X0 U465 ( .IN1(n438), .IN2(n434), .QN(n442) );
  XOR2X1 U466 ( .IN1(n443), .IN2(G13), .Q(G1336) );
  NAND2X0 U467 ( .IN1(n438), .IN2(n444), .QN(n443) );
  AND3X1 U468 ( .IN1(n419), .IN2(n411), .IN3(n445), .Q(n438) );
  XOR2X1 U469 ( .IN1(n446), .IN2(G12), .Q(G1335) );
  NAND2X0 U470 ( .IN1(n447), .IN2(n439), .QN(n446) );
  XOR2X1 U471 ( .IN1(n448), .IN2(G11), .Q(G1334) );
  NAND2X0 U472 ( .IN1(n447), .IN2(n441), .QN(n448) );
  XOR2X1 U473 ( .IN1(n449), .IN2(G10), .Q(G1333) );
  NAND2X0 U474 ( .IN1(n447), .IN2(n434), .QN(n449) );
  XOR2X1 U475 ( .IN1(n450), .IN2(G9), .Q(G1332) );
  NAND2X0 U476 ( .IN1(n447), .IN2(n444), .QN(n450) );
  AND3X1 U477 ( .IN1(n421), .IN2(n451), .IN3(n445), .Q(n447) );
  AND3X1 U478 ( .IN1(n452), .IN2(n453), .IN3(n430), .Q(n445) );
  XNOR2X1 U479 ( .IN1(G8), .IN2(n454), .Q(G1331) );
  NOR2X0 U480 ( .IN1(n455), .IN2(n416), .QN(n454) );
  XNOR2X1 U481 ( .IN1(G7), .IN2(n456), .Q(G1330) );
  NOR2X0 U482 ( .IN1(n457), .IN2(n416), .QN(n456) );
  XNOR2X1 U483 ( .IN1(G6), .IN2(n458), .Q(G1329) );
  NOR2X0 U484 ( .IN1(n459), .IN2(n416), .QN(n458) );
  NAND4X0 U485 ( .IN1(n432), .IN2(n425), .IN3(n460), .IN4(n419), .QN(n416) );
  AND2X1 U486 ( .IN1(n453), .IN2(n411), .Q(n460) );
  XOR2X1 U487 ( .IN1(n461), .IN2(G3), .Q(G1326) );
  NAND2X0 U488 ( .IN1(n462), .IN2(n441), .QN(n461) );
  XOR2X1 U489 ( .IN1(n463), .IN2(G2), .Q(G1325) );
  NAND2X0 U490 ( .IN1(n462), .IN2(n434), .QN(n463) );
  XOR2X1 U491 ( .IN1(n464), .IN2(G1), .Q(G1324) );
  NAND2X0 U492 ( .IN1(n462), .IN2(n444), .QN(n464) );
  XOR3X1 U493 ( .IN1(keyinput127), .IN2(keyinput118), .IN3(n465), .Q(G1355) );
  NOR2X0 U494 ( .IN1(n466), .IN2(n467), .QN(n465) );
  XOR2X1 U495 ( .IN1(keyinput110), .IN2(n468), .Q(n467) );
  AND2X1 U496 ( .IN1(n469), .IN2(n470), .Q(n468) );
  XOR2X1 U497 ( .IN1(n471), .IN2(keyinput109), .Q(n466) );
  NAND2X0 U498 ( .IN1(G32), .IN2(n470), .QN(n471) );
  XNOR2X1 U499 ( .IN1(n472), .IN2(keyinput95), .Q(n470) );
  NAND2X0 U500 ( .IN1(G32), .IN2(n469), .QN(n472) );
  XNOR2X1 U501 ( .IN1(n473), .IN2(keyinput87), .Q(n469) );
  NAND2X0 U502 ( .IN1(n422), .IN2(n411), .QN(n473) );
  XOR2X1 U503 ( .IN1(keyinput117), .IN2(n474), .Q(G1352) );
  OA21X1 U504 ( .IN1(n475), .IN2(n476), .IN3(n477), .Q(n474) );
  XOR2X1 U505 ( .IN1(keyinput108), .IN2(n478), .Q(n477) );
  NOR2X0 U506 ( .IN1(n475), .IN2(n479), .QN(n478) );
  XOR2X1 U507 ( .IN1(n480), .IN2(keyinput94), .Q(n475) );
  OR2X1 U508 ( .IN1(n476), .IN2(n479), .Q(n480) );
  INVX0 U509 ( .INP(G29), .ZN(n479) );
  XNOR2X1 U510 ( .IN1(n481), .IN2(keyinput86), .Q(n476) );
  NAND2X0 U511 ( .IN1(n422), .IN2(n432), .QN(n481) );
  INVX0 U512 ( .INP(n420), .ZN(n422) );
  XOR2X1 U513 ( .IN1(n482), .IN2(keyinput79), .Q(n420) );
  NAND3X0 U514 ( .IN1(n434), .IN2(n415), .IN3(n483), .QN(n482) );
  XOR3X1 U515 ( .IN1(keyinput126), .IN2(keyinput116), .IN3(n484), .Q(G1347) );
  NAND2X0 U516 ( .IN1(n485), .IN2(n486), .QN(n484) );
  XOR2X1 U517 ( .IN1(keyinput106), .IN2(n487), .Q(n486) );
  NOR2X0 U518 ( .IN1(n488), .IN2(n489), .QN(n487) );
  XOR2X1 U519 ( .IN1(keyinput107), .IN2(n490), .Q(n485) );
  NOR2X0 U520 ( .IN1(n488), .IN2(n491), .QN(n490) );
  XOR2X1 U521 ( .IN1(n492), .IN2(keyinput93), .Q(n488) );
  OR2X1 U522 ( .IN1(n491), .IN2(n489), .Q(n492) );
  XNOR2X1 U523 ( .IN1(n493), .IN2(keyinput85), .Q(n491) );
  NAND2X0 U524 ( .IN1(n494), .IN2(n411), .QN(n493) );
  XOR3X1 U525 ( .IN1(keyinput125), .IN2(keyinput115), .IN3(n495), .Q(G1346) );
  NOR2X0 U526 ( .IN1(n496), .IN2(n497), .QN(n495) );
  XOR2X1 U527 ( .IN1(n498), .IN2(keyinput105), .Q(n497) );
  NAND2X0 U528 ( .IN1(n499), .IN2(n500), .QN(n498) );
  XOR2X1 U529 ( .IN1(n501), .IN2(keyinput104), .Q(n496) );
  NAND2X0 U530 ( .IN1(G23), .IN2(n499), .QN(n501) );
  XNOR2X1 U531 ( .IN1(n502), .IN2(keyinput92), .Q(n499) );
  NAND2X0 U532 ( .IN1(G23), .IN2(n500), .QN(n502) );
  XNOR2X1 U533 ( .IN1(n503), .IN2(keyinput84), .Q(n500) );
  NAND2X0 U534 ( .IN1(n421), .IN2(n494), .QN(n503) );
  XOR3X1 U535 ( .IN1(keyinput124), .IN2(keyinput114), .IN3(n504), .Q(G1345) );
  NAND2X0 U536 ( .IN1(n505), .IN2(n506), .QN(n504) );
  XOR2X1 U537 ( .IN1(keyinput102), .IN2(n507), .Q(n506) );
  NOR2X0 U538 ( .IN1(n508), .IN2(n509), .QN(n507) );
  XOR2X1 U539 ( .IN1(keyinput103), .IN2(n510), .Q(n505) );
  NOR2X0 U540 ( .IN1(n511), .IN2(n509), .QN(n510) );
  XNOR2X1 U541 ( .IN1(n512), .IN2(keyinput91), .Q(n509) );
  OR2X1 U542 ( .IN1(n511), .IN2(n508), .Q(n512) );
  XNOR2X1 U543 ( .IN1(n513), .IN2(keyinput83), .Q(n511) );
  NAND2X0 U544 ( .IN1(n430), .IN2(n494), .QN(n513) );
  XOR3X1 U545 ( .IN1(keyinput123), .IN2(keyinput113), .IN3(n514), .Q(G1344) );
  NAND2X0 U546 ( .IN1(n515), .IN2(n516), .QN(n514) );
  XOR2X1 U547 ( .IN1(keyinput100), .IN2(n517), .Q(n516) );
  AND2X1 U548 ( .IN1(G21), .IN2(n518), .Q(n517) );
  XOR2X1 U549 ( .IN1(n519), .IN2(keyinput101), .Q(n515) );
  NAND2X0 U550 ( .IN1(n518), .IN2(n520), .QN(n519) );
  XOR2X1 U551 ( .IN1(n521), .IN2(keyinput90), .Q(n518) );
  NAND2X0 U552 ( .IN1(n520), .IN2(G21), .QN(n521) );
  XOR2X1 U553 ( .IN1(n522), .IN2(keyinput82), .Q(n520) );
  NAND2X0 U554 ( .IN1(n494), .IN2(n432), .QN(n522) );
  XNOR2X1 U555 ( .IN1(n523), .IN2(keyinput78), .Q(n494) );
  NAND3X0 U556 ( .IN1(n444), .IN2(n459), .IN3(n483), .QN(n523) );
  AND3X1 U557 ( .IN1(n524), .IN2(n457), .IN3(n439), .Q(n483) );
  XOR3X1 U558 ( .IN1(keyinput121), .IN2(keyinput111), .IN3(n525), .Q(G1340) );
  NAND2X0 U559 ( .IN1(n526), .IN2(n527), .QN(n525) );
  XOR2X1 U560 ( .IN1(keyinput97), .IN2(n528), .Q(n527) );
  AND2X1 U561 ( .IN1(n529), .IN2(n530), .Q(n528) );
  XOR2X1 U562 ( .IN1(n531), .IN2(keyinput96), .Q(n526) );
  NAND2X0 U563 ( .IN1(G17), .IN2(n530), .QN(n531) );
  XNOR2X1 U564 ( .IN1(n532), .IN2(keyinput88), .Q(n530) );
  NAND2X0 U565 ( .IN1(G17), .IN2(n529), .QN(n532) );
  XNOR2X1 U566 ( .IN1(n533), .IN2(keyinput80), .Q(n529) );
  NAND2X0 U567 ( .IN1(n410), .IN2(n432), .QN(n533) );
  XOR2X1 U568 ( .IN1(n534), .IN2(keyinput77), .Q(n410) );
  NAND3X0 U569 ( .IN1(n444), .IN2(n459), .IN3(n433), .QN(n534) );
  AND3X1 U570 ( .IN1(n441), .IN2(n455), .IN3(n524), .Q(n433) );
  XOR2X1 U571 ( .IN1(n535), .IN2(keyinput76), .Q(n524) );
  NAND3X0 U572 ( .IN1(n536), .IN2(n537), .IN3(n538), .QN(n535) );
  OA222X1 U573 ( .IN1(n539), .IN2(n540), .IN3(n541), .IN4(n542), .IN5(n543), 
        .IN6(n430), .Q(n538) );
  OA22X1 U574 ( .IN1(n411), .IN2(n544), .IN3(keyinput72), .IN4(n545), .Q(n543)
         );
  MUX21X1 U575 ( .IN1(n546), .IN2(n547), .S(n419), .Q(n544) );
  NAND2X0 U576 ( .IN1(keyinput71), .IN2(keyinput75), .QN(n547) );
  OA22X1 U577 ( .IN1(n548), .IN2(n549), .IN3(keyinput73), .IN4(n550), .Q(n546)
         );
  OR2X1 U578 ( .IN1(n452), .IN2(keyinput71), .Q(n549) );
  INVX0 U579 ( .INP(keyinput72), .ZN(n542) );
  NOR2X0 U580 ( .IN1(n430), .IN2(n545), .QN(n541) );
  NAND3X0 U581 ( .IN1(n551), .IN2(n411), .IN3(n552), .QN(n545) );
  XOR2X1 U582 ( .IN1(keyinput66), .IN2(n432), .Q(n552) );
  INVX0 U583 ( .INP(n451), .ZN(n411) );
  XOR2X1 U584 ( .IN1(keyinput67), .IN2(n419), .Q(n551) );
  INVX0 U585 ( .INP(n421), .ZN(n419) );
  INVX0 U586 ( .INP(keyinput73), .ZN(n540) );
  NOR2X0 U587 ( .IN1(n553), .IN2(n550), .QN(n539) );
  XOR2X1 U588 ( .IN1(keyinput68), .IN2(n432), .Q(n550) );
  NAND2X0 U589 ( .IN1(n554), .IN2(n548), .QN(n537) );
  INVX0 U590 ( .INP(keyinput75), .ZN(n548) );
  NAND4X0 U591 ( .IN1(n555), .IN2(n451), .IN3(n432), .IN4(n425), .QN(n554) );
  XOR2X1 U592 ( .IN1(n421), .IN2(keyinput71), .Q(n555) );
  XOR2X1 U593 ( .IN1(n556), .IN2(keyinput74), .Q(n536) );
  NAND4X0 U594 ( .IN1(n430), .IN2(n557), .IN3(n451), .IN4(n558), .QN(n556) );
  XOR2X1 U595 ( .IN1(keyinput69), .IN2(n432), .Q(n558) );
  XOR2X1 U596 ( .IN1(n421), .IN2(keyinput70), .Q(n557) );
  XOR2X1 U597 ( .IN1(n559), .IN2(keyinput119), .Q(G1327) );
  MUX21X1 U598 ( .IN1(n560), .IN2(n561), .S(G4), .Q(n559) );
  NOR2X0 U599 ( .IN1(n455), .IN2(n562), .QN(n561) );
  NAND2X0 U600 ( .IN1(n462), .IN2(n439), .QN(n560) );
  INVX0 U601 ( .INP(n562), .ZN(n462) );
  NAND3X0 U602 ( .IN1(n432), .IN2(n453), .IN3(n563), .QN(n562) );
  INVX0 U603 ( .INP(n553), .ZN(n563) );
  NAND3X0 U604 ( .IN1(n421), .IN2(n425), .IN3(n451), .QN(n553) );
  XOR2X1 U605 ( .IN1(n564), .IN2(n565), .Q(n451) );
  XOR3X1 U606 ( .IN1(G24), .IN2(G20), .IN3(n566), .Q(n565) );
  OA21X1 U607 ( .IN1(n567), .IN2(n568), .IN3(n569), .Q(n566) );
  NAND3X0 U608 ( .IN1(G40), .IN2(n568), .IN3(G41), .QN(n569) );
  XNOR2X1 U609 ( .IN1(n570), .IN2(n571), .Q(n568) );
  AND2X1 U610 ( .IN1(G40), .IN2(G41), .Q(n567) );
  XNOR3X1 U611 ( .IN1(keyinput62), .IN2(G32), .IN3(G28), .Q(n564) );
  INVX0 U612 ( .INP(n430), .ZN(n425) );
  MUX21X1 U613 ( .IN1(n572), .IN2(n573), .S(n574), .Q(n430) );
  XOR3X1 U614 ( .IN1(G22), .IN2(G18), .IN3(n575), .Q(n574) );
  XOR2X1 U615 ( .IN1(G30), .IN2(G26), .Q(n575) );
  NAND2X0 U616 ( .IN1(n576), .IN2(n577), .QN(n573) );
  AND2X1 U617 ( .IN1(n577), .IN2(n576), .Q(n572) );
  NAND3X0 U618 ( .IN1(G41), .IN2(n578), .IN3(G38), .QN(n576) );
  AO21X1 U619 ( .IN1(G38), .IN2(G41), .IN3(n578), .Q(n577) );
  XNOR2X1 U620 ( .IN1(n571), .IN2(n579), .Q(n578) );
  XOR3X1 U621 ( .IN1(G14), .IN2(G13), .IN3(n580), .Q(n571) );
  XOR2X1 U622 ( .IN1(n581), .IN2(G16), .Q(n580) );
  INVX0 U623 ( .INP(G15), .ZN(n581) );
  XOR2X1 U624 ( .IN1(n582), .IN2(keyinput63), .Q(n421) );
  NAND2X0 U625 ( .IN1(n583), .IN2(n584), .QN(n582) );
  XOR2X1 U626 ( .IN1(n585), .IN2(keyinput61), .Q(n584) );
  NAND2X0 U627 ( .IN1(n586), .IN2(n587), .QN(n585) );
  XOR2X1 U628 ( .IN1(n588), .IN2(keyinput60), .Q(n583) );
  NAND2X0 U629 ( .IN1(n586), .IN2(n589), .QN(n588) );
  XOR2X1 U630 ( .IN1(n590), .IN2(keyinput57), .Q(n586) );
  NAND2X0 U631 ( .IN1(n587), .IN2(n589), .QN(n590) );
  XNOR3X1 U632 ( .IN1(G23), .IN2(G19), .IN3(n591), .Q(n589) );
  XNOR2X1 U633 ( .IN1(G27), .IN2(G31), .Q(n591) );
  XOR2X1 U634 ( .IN1(n592), .IN2(keyinput55), .Q(n587) );
  NAND2X0 U635 ( .IN1(n593), .IN2(n594), .QN(n592) );
  XOR2X1 U636 ( .IN1(keyinput52), .IN2(n595), .Q(n594) );
  NOR2X0 U637 ( .IN1(n596), .IN2(n597), .QN(n595) );
  XOR2X1 U638 ( .IN1(keyinput49), .IN2(n598), .Q(n597) );
  XOR2X1 U639 ( .IN1(n599), .IN2(keyinput53), .Q(n593) );
  NAND2X0 U640 ( .IN1(n600), .IN2(n601), .QN(n599) );
  INVX0 U641 ( .INP(n602), .ZN(n601) );
  XNOR2X1 U642 ( .IN1(keyinput49), .IN2(n598), .Q(n600) );
  NOR2X0 U643 ( .IN1(n596), .IN2(n602), .QN(n598) );
  XOR2X1 U644 ( .IN1(n603), .IN2(keyinput47), .Q(n602) );
  NAND2X0 U645 ( .IN1(n604), .IN2(n605), .QN(n603) );
  XOR2X1 U646 ( .IN1(n606), .IN2(keyinput44), .Q(n605) );
  NAND2X0 U647 ( .IN1(n607), .IN2(n608), .QN(n606) );
  XOR2X1 U648 ( .IN1(n609), .IN2(keyinput45), .Q(n604) );
  NAND2X0 U649 ( .IN1(n607), .IN2(n579), .QN(n609) );
  XOR2X1 U650 ( .IN1(n610), .IN2(keyinput41), .Q(n607) );
  NAND2X0 U651 ( .IN1(n608), .IN2(n579), .QN(n610) );
  XNOR2X1 U652 ( .IN1(n611), .IN2(keyinput38), .Q(n579) );
  NAND2X0 U653 ( .IN1(n612), .IN2(n613), .QN(n611) );
  XOR2X1 U654 ( .IN1(keyinput34), .IN2(n614), .Q(n613) );
  NOR2X0 U655 ( .IN1(n615), .IN2(n616), .QN(n614) );
  XNOR2X1 U656 ( .IN1(keyinput24), .IN2(n617), .Q(n615) );
  XOR2X1 U657 ( .IN1(keyinput35), .IN2(n618), .Q(n612) );
  NOR2X0 U658 ( .IN1(n619), .IN2(n616), .QN(n618) );
  XNOR2X1 U659 ( .IN1(n620), .IN2(keyinput29), .Q(n616) );
  NAND2X0 U660 ( .IN1(n621), .IN2(n622), .QN(n620) );
  XOR2X1 U661 ( .IN1(keyinput24), .IN2(n617), .Q(n622) );
  AND2X1 U662 ( .IN1(n623), .IN2(n624), .Q(n617) );
  XOR2X1 U663 ( .IN1(n625), .IN2(keyinput15), .Q(n624) );
  NAND2X0 U664 ( .IN1(G9), .IN2(n626), .QN(n625) );
  XOR2X1 U665 ( .IN1(n627), .IN2(keyinput16), .Q(n623) );
  NAND2X0 U666 ( .IN1(G10), .IN2(n626), .QN(n627) );
  XNOR2X1 U667 ( .IN1(n628), .IN2(keyinput5), .Q(n626) );
  NAND2X0 U668 ( .IN1(G9), .IN2(G10), .QN(n628) );
  XOR2X1 U669 ( .IN1(keyinput25), .IN2(n629), .Q(n621) );
  XNOR2X1 U670 ( .IN1(keyinput25), .IN2(n629), .Q(n619) );
  AND2X1 U671 ( .IN1(n630), .IN2(n631), .Q(n629) );
  XOR2X1 U672 ( .IN1(keyinput17), .IN2(n632), .Q(n631) );
  NOR2X0 U673 ( .IN1(n633), .IN2(n634), .QN(n632) );
  INVX0 U674 ( .INP(G11), .ZN(n633) );
  XOR2X1 U675 ( .IN1(keyinput18), .IN2(n635), .Q(n630) );
  NOR2X0 U676 ( .IN1(n636), .IN2(n634), .QN(n635) );
  XNOR2X1 U677 ( .IN1(n637), .IN2(keyinput6), .Q(n634) );
  NAND2X0 U678 ( .IN1(G11), .IN2(G12), .QN(n637) );
  INVX0 U679 ( .INP(G12), .ZN(n636) );
  XNOR2X1 U680 ( .IN1(n638), .IN2(keyinput0), .Q(n596) );
  NAND2X0 U681 ( .IN1(G39), .IN2(G41), .QN(n638) );
  NAND2X0 U682 ( .IN1(n639), .IN2(n640), .QN(n453) );
  NAND3X0 U683 ( .IN1(n457), .IN2(n455), .IN3(n641), .QN(n640) );
  NAND2X0 U684 ( .IN1(n434), .IN2(n444), .QN(n641) );
  INVX0 U685 ( .INP(n441), .ZN(n457) );
  NAND3X0 U686 ( .IN1(n459), .IN2(n415), .IN3(n642), .QN(n639) );
  XOR2X1 U687 ( .IN1(n643), .IN2(n455), .Q(n642) );
  INVX0 U688 ( .INP(n439), .ZN(n455) );
  MUX21X1 U689 ( .IN1(n644), .IN2(n645), .S(n646), .Q(n439) );
  XOR3X1 U690 ( .IN1(G16), .IN2(G12), .IN3(n647), .Q(n646) );
  XOR2X1 U691 ( .IN1(G8), .IN2(G4), .Q(n647) );
  NAND2X0 U692 ( .IN1(n648), .IN2(n649), .QN(n645) );
  AND2X1 U693 ( .IN1(n649), .IN2(n648), .Q(n644) );
  NAND3X0 U694 ( .IN1(G41), .IN2(n650), .IN3(G36), .QN(n648) );
  AO21X1 U695 ( .IN1(G36), .IN2(G41), .IN3(n650), .Q(n649) );
  XOR2X1 U696 ( .IN1(n651), .IN2(n652), .Q(n650) );
  NAND2X0 U697 ( .IN1(keyinput65), .IN2(n441), .QN(n643) );
  MUX21X1 U698 ( .IN1(n653), .IN2(n654), .S(n655), .Q(n441) );
  XOR3X1 U699 ( .IN1(G15), .IN2(G11), .IN3(n656), .Q(n655) );
  XOR2X1 U700 ( .IN1(G7), .IN2(G3), .Q(n656) );
  NAND2X0 U701 ( .IN1(n657), .IN2(n658), .QN(n654) );
  AND2X1 U702 ( .IN1(n658), .IN2(n657), .Q(n653) );
  NAND3X0 U703 ( .IN1(G41), .IN2(n659), .IN3(G35), .QN(n657) );
  AO21X1 U704 ( .IN1(G35), .IN2(G41), .IN3(n659), .Q(n658) );
  XOR2X1 U705 ( .IN1(n660), .IN2(n661), .Q(n659) );
  INVX0 U706 ( .INP(n444), .ZN(n415) );
  MUX21X1 U707 ( .IN1(n662), .IN2(n663), .S(n664), .Q(n444) );
  XOR3X1 U708 ( .IN1(G13), .IN2(G1), .IN3(n665), .Q(n664) );
  XOR2X1 U709 ( .IN1(G9), .IN2(G5), .Q(n665) );
  NAND2X0 U710 ( .IN1(n666), .IN2(n667), .QN(n663) );
  AND2X1 U711 ( .IN1(n667), .IN2(n666), .Q(n662) );
  NAND3X0 U712 ( .IN1(G41), .IN2(n668), .IN3(G33), .QN(n666) );
  AO21X1 U713 ( .IN1(G33), .IN2(G41), .IN3(n668), .Q(n667) );
  XOR2X1 U714 ( .IN1(n661), .IN2(n652), .Q(n668) );
  XOR3X1 U715 ( .IN1(n508), .IN2(G21), .IN3(n669), .Q(n652) );
  XOR2X1 U716 ( .IN1(G23), .IN2(n489), .Q(n669) );
  INVX0 U717 ( .INP(G24), .ZN(n489) );
  INVX0 U718 ( .INP(G22), .ZN(n508) );
  XNOR3X1 U719 ( .IN1(G18), .IN2(G17), .IN3(n670), .Q(n661) );
  XNOR2X1 U720 ( .IN1(G19), .IN2(G20), .Q(n670) );
  INVX0 U721 ( .INP(n434), .ZN(n459) );
  MUX21X1 U722 ( .IN1(n671), .IN2(n672), .S(n673), .Q(n434) );
  XOR3X1 U723 ( .IN1(G14), .IN2(G10), .IN3(n674), .Q(n673) );
  XOR2X1 U724 ( .IN1(G6), .IN2(G2), .Q(n674) );
  NAND2X0 U725 ( .IN1(n675), .IN2(n676), .QN(n672) );
  AND2X1 U726 ( .IN1(n676), .IN2(n675), .Q(n671) );
  NAND3X0 U727 ( .IN1(G41), .IN2(n677), .IN3(G34), .QN(n675) );
  AO21X1 U728 ( .IN1(G34), .IN2(G41), .IN3(n677), .Q(n676) );
  XOR2X1 U729 ( .IN1(n660), .IN2(n651), .Q(n677) );
  XOR3X1 U730 ( .IN1(n423), .IN2(G29), .IN3(n678), .Q(n651) );
  XNOR3X1 U731 ( .IN1(keyinput26), .IN2(G32), .IN3(G31), .Q(n678) );
  INVX0 U732 ( .INP(G30), .ZN(n423) );
  XOR3X1 U733 ( .IN1(G26), .IN2(n679), .IN3(n680), .Q(n660) );
  XNOR2X1 U734 ( .IN1(G27), .IN2(G28), .Q(n680) );
  INVX0 U735 ( .INP(n452), .ZN(n432) );
  XOR2X1 U736 ( .IN1(n681), .IN2(keyinput64), .Q(n452) );
  NAND2X0 U737 ( .IN1(n682), .IN2(n683), .QN(n681) );
  XOR2X1 U738 ( .IN1(keyinput59), .IN2(n684), .Q(n683) );
  NOR2X0 U739 ( .IN1(n685), .IN2(n686), .QN(n684) );
  XNOR2X1 U740 ( .IN1(keyinput54), .IN2(n687), .Q(n686) );
  INVX0 U741 ( .INP(n688), .ZN(n685) );
  XOR2X1 U742 ( .IN1(n689), .IN2(keyinput58), .Q(n682) );
  NAND2X0 U743 ( .IN1(n688), .IN2(n690), .QN(n689) );
  XOR2X1 U744 ( .IN1(n691), .IN2(keyinput56), .Q(n688) );
  NAND2X0 U745 ( .IN1(n692), .IN2(n690), .QN(n691) );
  XOR3X1 U746 ( .IN1(keyinput39), .IN2(G21), .IN3(n693), .Q(n690) );
  XNOR2X1 U747 ( .IN1(G17), .IN2(n694), .Q(n693) );
  OA21X1 U748 ( .IN1(G29), .IN2(n679), .IN3(n695), .Q(n694) );
  XOR2X1 U749 ( .IN1(n696), .IN2(keyinput19), .Q(n695) );
  NAND2X0 U750 ( .IN1(G29), .IN2(n679), .QN(n696) );
  INVX0 U751 ( .INP(G25), .ZN(n679) );
  XOR2X1 U752 ( .IN1(n687), .IN2(keyinput54), .Q(n692) );
  NAND2X0 U753 ( .IN1(n697), .IN2(n698), .QN(n687) );
  XOR2X1 U754 ( .IN1(keyinput50), .IN2(n699), .Q(n698) );
  NOR2X0 U755 ( .IN1(n700), .IN2(n701), .QN(n699) );
  XOR2X1 U756 ( .IN1(keyinput51), .IN2(n702), .Q(n697) );
  NOR2X0 U757 ( .IN1(n700), .IN2(n703), .QN(n702) );
  XNOR2X1 U758 ( .IN1(keyinput46), .IN2(n704), .Q(n703) );
  XOR2X1 U759 ( .IN1(n705), .IN2(keyinput48), .Q(n700) );
  NAND2X0 U760 ( .IN1(n706), .IN2(n707), .QN(n705) );
  INVX0 U761 ( .INP(n701), .ZN(n707) );
  NAND2X0 U762 ( .IN1(G37), .IN2(G41), .QN(n701) );
  XOR2X1 U763 ( .IN1(n704), .IN2(keyinput46), .Q(n706) );
  NAND2X0 U764 ( .IN1(n708), .IN2(n709), .QN(n704) );
  XOR2X1 U765 ( .IN1(n710), .IN2(keyinput42), .Q(n709) );
  NAND2X0 U766 ( .IN1(n711), .IN2(n608), .QN(n710) );
  XOR2X1 U767 ( .IN1(n712), .IN2(keyinput43), .Q(n708) );
  NAND2X0 U768 ( .IN1(n711), .IN2(n570), .QN(n712) );
  XOR2X1 U769 ( .IN1(n713), .IN2(keyinput40), .Q(n711) );
  NAND2X0 U770 ( .IN1(n608), .IN2(n570), .QN(n713) );
  XNOR2X1 U771 ( .IN1(n714), .IN2(keyinput37), .Q(n570) );
  NAND2X0 U772 ( .IN1(n715), .IN2(n716), .QN(n714) );
  XOR2X1 U773 ( .IN1(keyinput33), .IN2(n717), .Q(n716) );
  NOR2X0 U774 ( .IN1(n718), .IN2(n719), .QN(n717) );
  XOR2X1 U775 ( .IN1(n720), .IN2(keyinput23), .Q(n719) );
  XOR2X1 U776 ( .IN1(n721), .IN2(keyinput32), .Q(n715) );
  NAND2X0 U777 ( .IN1(n722), .IN2(n723), .QN(n721) );
  INVX0 U778 ( .INP(n718), .ZN(n722) );
  XOR2X1 U779 ( .IN1(n724), .IN2(keyinput28), .Q(n718) );
  NAND2X0 U780 ( .IN1(n725), .IN2(n723), .QN(n724) );
  XNOR2X1 U781 ( .IN1(n726), .IN2(keyinput22), .Q(n723) );
  NAND2X0 U782 ( .IN1(n727), .IN2(n728), .QN(n726) );
  XOR2X1 U783 ( .IN1(n729), .IN2(keyinput11), .Q(n728) );
  NAND2X0 U784 ( .IN1(G5), .IN2(n730), .QN(n729) );
  XOR2X1 U785 ( .IN1(n731), .IN2(keyinput12), .Q(n727) );
  NAND2X0 U786 ( .IN1(G6), .IN2(n730), .QN(n731) );
  XNOR2X1 U787 ( .IN1(n732), .IN2(keyinput3), .Q(n730) );
  NAND2X0 U788 ( .IN1(G6), .IN2(G5), .QN(n732) );
  XNOR2X1 U789 ( .IN1(keyinput23), .IN2(n720), .Q(n725) );
  NAND2X0 U790 ( .IN1(n733), .IN2(n734), .QN(n720) );
  XOR2X1 U791 ( .IN1(keyinput14), .IN2(n735), .Q(n734) );
  AND2X1 U792 ( .IN1(n736), .IN2(G8), .Q(n735) );
  XOR2X1 U793 ( .IN1(n737), .IN2(keyinput13), .Q(n733) );
  NAND2X0 U794 ( .IN1(G7), .IN2(n736), .QN(n737) );
  XNOR2X1 U795 ( .IN1(n738), .IN2(keyinput4), .Q(n736) );
  NAND2X0 U796 ( .IN1(G8), .IN2(G7), .QN(n738) );
  XOR2X1 U797 ( .IN1(n739), .IN2(keyinput36), .Q(n608) );
  NAND2X0 U798 ( .IN1(n740), .IN2(n741), .QN(n739) );
  XOR2X1 U799 ( .IN1(n742), .IN2(keyinput31), .Q(n741) );
  NAND2X0 U800 ( .IN1(n743), .IN2(n744), .QN(n742) );
  XOR2X1 U801 ( .IN1(n745), .IN2(keyinput30), .Q(n740) );
  NAND2X0 U802 ( .IN1(n746), .IN2(n744), .QN(n745) );
  XNOR2X1 U803 ( .IN1(n747), .IN2(keyinput27), .Q(n744) );
  NAND2X0 U804 ( .IN1(n743), .IN2(n746), .QN(n747) );
  XOR2X1 U805 ( .IN1(n748), .IN2(keyinput21), .Q(n743) );
  NAND2X0 U806 ( .IN1(n749), .IN2(n750), .QN(n748) );
  XOR2X1 U807 ( .IN1(keyinput10), .IN2(n751), .Q(n750) );
  AND2X1 U808 ( .IN1(G4), .IN2(n752), .Q(n751) );
  XOR2X1 U809 ( .IN1(n753), .IN2(keyinput9), .Q(n749) );
  NAND2X0 U810 ( .IN1(n752), .IN2(G3), .QN(n753) );
  XOR2X1 U811 ( .IN1(n754), .IN2(keyinput2), .Q(n752) );
  NAND2X0 U812 ( .IN1(G3), .IN2(G4), .QN(n754) );
  XOR2X1 U813 ( .IN1(n755), .IN2(keyinput20), .Q(n746) );
  NAND2X0 U814 ( .IN1(n756), .IN2(n757), .QN(n755) );
  XOR2X1 U815 ( .IN1(n758), .IN2(keyinput7), .Q(n757) );
  NAND2X0 U816 ( .IN1(n759), .IN2(G1), .QN(n758) );
  XOR2X1 U817 ( .IN1(n760), .IN2(keyinput8), .Q(n756) );
  NAND2X0 U818 ( .IN1(n759), .IN2(G2), .QN(n760) );
  XOR2X1 U819 ( .IN1(n761), .IN2(keyinput1), .Q(n759) );
  NAND2X0 U820 ( .IN1(G2), .IN2(G1), .QN(n761) );
endmodule

