
module c499 ( N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, 
        N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, 
        N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, 
        N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, 
        N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, 
        N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, keyinput0, 
        keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, 
        keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, 
        keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, 
        keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, 
        keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, 
        keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, 
        keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, 
        keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, 
        keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, 
        keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, 
        keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, 
        keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, 
        keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, 
        keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, 
        keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, 
        keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, 
        keyinput97, keyinput98, keyinput99, keyinput100, keyinput101, 
        keyinput102, keyinput103, keyinput104, keyinput105, keyinput106, 
        keyinput107, keyinput108, keyinput109, keyinput110, keyinput111, 
        keyinput112, keyinput113, keyinput114, keyinput115, keyinput116, 
        keyinput117, keyinput118, keyinput119, keyinput120, keyinput121, 
        keyinput122, keyinput123, keyinput124, keyinput125, keyinput126, 
        keyinput127 );
  input N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57,
         N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109,
         N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135,
         N136, N137, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4,
         keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10,
         keyinput11, keyinput12, keyinput13, keyinput14, keyinput15,
         keyinput16, keyinput17, keyinput18, keyinput19, keyinput20,
         keyinput21, keyinput22, keyinput23, keyinput24, keyinput25,
         keyinput26, keyinput27, keyinput28, keyinput29, keyinput30,
         keyinput31, keyinput32, keyinput33, keyinput34, keyinput35,
         keyinput36, keyinput37, keyinput38, keyinput39, keyinput40,
         keyinput41, keyinput42, keyinput43, keyinput44, keyinput45,
         keyinput46, keyinput47, keyinput48, keyinput49, keyinput50,
         keyinput51, keyinput52, keyinput53, keyinput54, keyinput55,
         keyinput56, keyinput57, keyinput58, keyinput59, keyinput60,
         keyinput61, keyinput62, keyinput63, keyinput64, keyinput65,
         keyinput66, keyinput67, keyinput68, keyinput69, keyinput70,
         keyinput71, keyinput72, keyinput73, keyinput74, keyinput75,
         keyinput76, keyinput77, keyinput78, keyinput79, keyinput80,
         keyinput81, keyinput82, keyinput83, keyinput84, keyinput85,
         keyinput86, keyinput87, keyinput88, keyinput89, keyinput90,
         keyinput91, keyinput92, keyinput93, keyinput94, keyinput95,
         keyinput96, keyinput97, keyinput98, keyinput99, keyinput100,
         keyinput101, keyinput102, keyinput103, keyinput104, keyinput105,
         keyinput106, keyinput107, keyinput108, keyinput109, keyinput110,
         keyinput111, keyinput112, keyinput113, keyinput114, keyinput115,
         keyinput116, keyinput117, keyinput118, keyinput119, keyinput120,
         keyinput121, keyinput122, keyinput123, keyinput124, keyinput125,
         keyinput126, keyinput127;
  output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745,
         N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
  wire   n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449;

  XOR3X1 U247 ( .IN1(keyinput126), .IN2(N121), .IN3(n227), .Q(N754) );
  NOR2X0 U248 ( .IN1(n228), .IN2(n229), .QN(n227) );
  XOR3X1 U249 ( .IN1(keyinput127), .IN2(N125), .IN3(n230), .Q(N755) );
  NOR2X0 U250 ( .IN1(n229), .IN2(n231), .QN(n230) );
  XOR3X1 U251 ( .IN1(n232), .IN2(n233), .IN3(n234), .Q(N753) );
  NAND2X0 U252 ( .IN1(n235), .IN2(n236), .QN(n234) );
  XOR2X1 U253 ( .IN1(keyinput125), .IN2(keyinput106), .Q(n232) );
  XOR3X1 U254 ( .IN1(n237), .IN2(n238), .IN3(n239), .Q(N752) );
  NAND2X0 U255 ( .IN1(n240), .IN2(n236), .QN(n239) );
  INVX0 U256 ( .INP(n229), .ZN(n236) );
  XOR2X1 U257 ( .IN1(n241), .IN2(keyinput85), .Q(n229) );
  NAND4X0 U258 ( .IN1(n242), .IN2(n243), .IN3(n244), .IN4(n245), .QN(n241) );
  XOR2X1 U259 ( .IN1(keyinput71), .IN2(n246), .Q(n244) );
  XOR2X1 U260 ( .IN1(keyinput124), .IN2(keyinput105), .Q(n237) );
  XOR2X1 U261 ( .IN1(n247), .IN2(n248), .Q(N751) );
  NAND2X0 U262 ( .IN1(n249), .IN2(n250), .QN(n248) );
  XOR3X1 U263 ( .IN1(N105), .IN2(n251), .IN3(n252), .Q(N750) );
  NAND2X0 U264 ( .IN1(n249), .IN2(n253), .QN(n252) );
  XOR2X1 U265 ( .IN1(keyinput123), .IN2(keyinput104), .Q(n251) );
  XOR3X1 U266 ( .IN1(keyinput103), .IN2(n254), .IN3(n255), .Q(N749) );
  NAND2X0 U267 ( .IN1(n249), .IN2(n235), .QN(n255) );
  XOR3X1 U268 ( .IN1(keyinput102), .IN2(n256), .IN3(n257), .Q(N748) );
  NAND2X0 U269 ( .IN1(n249), .IN2(n240), .QN(n257) );
  XOR2X1 U270 ( .IN1(n258), .IN2(keyinput84), .Q(n249) );
  NAND4X0 U271 ( .IN1(n243), .IN2(n246), .IN3(n245), .IN4(n259), .QN(n258) );
  XOR3X1 U272 ( .IN1(keyinput101), .IN2(N93), .IN3(n260), .Q(N747) );
  AND2X1 U273 ( .IN1(n261), .IN2(n250), .Q(n260) );
  XOR3X1 U274 ( .IN1(N89), .IN2(n262), .IN3(n263), .Q(N746) );
  NAND2X0 U275 ( .IN1(n261), .IN2(n253), .QN(n263) );
  XOR2X1 U276 ( .IN1(keyinput122), .IN2(keyinput100), .Q(n262) );
  XOR3X1 U277 ( .IN1(keyinput121), .IN2(N85), .IN3(n264), .Q(N745) );
  NAND2X0 U278 ( .IN1(n235), .IN2(n261), .QN(n264) );
  XOR3X1 U279 ( .IN1(N81), .IN2(n265), .IN3(n266), .Q(N744) );
  NAND2X0 U280 ( .IN1(n240), .IN2(n261), .QN(n266) );
  XNOR2X1 U281 ( .IN1(n267), .IN2(keyinput83), .Q(n261) );
  NAND4X0 U282 ( .IN1(n245), .IN2(n268), .IN3(n242), .IN4(n269), .QN(n267) );
  NOR2X0 U283 ( .IN1(n270), .IN2(n271), .QN(n269) );
  XOR2X1 U284 ( .IN1(keyinput70), .IN2(n246), .Q(n271) );
  XOR2X1 U285 ( .IN1(keyinput69), .IN2(n272), .Q(n270) );
  XOR2X1 U286 ( .IN1(keyinput99), .IN2(keyinput120), .Q(n265) );
  XNOR3X1 U287 ( .IN1(keyinput119), .IN2(N77), .IN3(n273), .Q(N743) );
  NAND2X0 U288 ( .IN1(n274), .IN2(n250), .QN(n273) );
  XOR3X1 U289 ( .IN1(keyinput98), .IN2(n275), .IN3(n276), .Q(N742) );
  NAND2X0 U290 ( .IN1(n274), .IN2(n253), .QN(n276) );
  XOR3X1 U291 ( .IN1(n277), .IN2(n278), .IN3(n279), .Q(N741) );
  NAND2X0 U292 ( .IN1(n274), .IN2(n235), .QN(n279) );
  XOR2X1 U293 ( .IN1(keyinput97), .IN2(keyinput118), .Q(n277) );
  XOR3X1 U294 ( .IN1(N65), .IN2(n280), .IN3(n281), .Q(N740) );
  NAND2X0 U295 ( .IN1(n274), .IN2(n240), .QN(n281) );
  XOR2X1 U296 ( .IN1(n282), .IN2(keyinput82), .Q(n274) );
  NAND4X0 U297 ( .IN1(n245), .IN2(n268), .IN3(n246), .IN4(n283), .QN(n282) );
  NOR2X0 U298 ( .IN1(n284), .IN2(n285), .QN(n283) );
  XOR2X1 U299 ( .IN1(keyinput68), .IN2(n259), .Q(n285) );
  XOR2X1 U300 ( .IN1(keyinput67), .IN2(n272), .Q(n284) );
  XNOR2X1 U301 ( .IN1(n286), .IN2(keyinput79), .Q(n245) );
  AO221X1 U302 ( .IN1(n287), .IN2(n288), .IN3(n289), .IN4(n290), .IN5(n291), 
        .Q(n286) );
  MUX21X1 U303 ( .IN1(n292), .IN2(n293), .S(n294), .Q(n291) );
  NAND4X0 U304 ( .IN1(keyinput77), .IN2(n295), .IN3(n296), .IN4(n297), .QN(
        n293) );
  NAND3X0 U305 ( .IN1(n298), .IN2(n253), .IN3(n299), .QN(n297) );
  XOR2X1 U306 ( .IN1(n250), .IN2(keyinput61), .Q(n299) );
  NAND2X0 U307 ( .IN1(keyinput62), .IN2(n300), .QN(n296) );
  INVX0 U308 ( .INP(n301), .ZN(n300) );
  OR2X1 U309 ( .IN1(n287), .IN2(n288), .Q(n295) );
  OAI221X1 U310 ( .IN1(n301), .IN2(keyinput62), .IN3(n290), .IN4(n289), .IN5(
        keyinput76), .QN(n292) );
  NAND3X0 U311 ( .IN1(n235), .IN2(n302), .IN3(n303), .QN(n301) );
  XOR2X1 U312 ( .IN1(n250), .IN2(keyinput64), .Q(n303) );
  XOR2X1 U313 ( .IN1(keyinput63), .IN2(n253), .Q(n302) );
  INVX0 U314 ( .INP(keyinput77), .ZN(n290) );
  NAND3X0 U315 ( .IN1(n304), .IN2(n298), .IN3(n305), .QN(n289) );
  XOR2X1 U316 ( .IN1(n228), .IN2(keyinput65), .Q(n305) );
  XOR2X1 U317 ( .IN1(keyinput66), .IN2(n231), .Q(n304) );
  INVX0 U318 ( .INP(keyinput76), .ZN(n288) );
  NAND3X0 U319 ( .IN1(n250), .IN2(n306), .IN3(n307), .QN(n287) );
  XOR2X1 U320 ( .IN1(n228), .IN2(keyinput60), .Q(n307) );
  XOR2X1 U321 ( .IN1(keyinput59), .IN2(n298), .Q(n306) );
  XOR2X1 U322 ( .IN1(keyinput96), .IN2(keyinput117), .Q(n280) );
  XOR3X1 U323 ( .IN1(N61), .IN2(n308), .IN3(n309), .Q(N739) );
  NAND2X0 U324 ( .IN1(n310), .IN2(n242), .QN(n309) );
  XOR2X1 U325 ( .IN1(keyinput95), .IN2(keyinput116), .Q(n308) );
  XNOR3X1 U326 ( .IN1(n311), .IN2(N57), .IN3(n312), .Q(N738) );
  NAND2X0 U327 ( .IN1(n310), .IN2(n246), .QN(n312) );
  XOR2X1 U328 ( .IN1(keyinput94), .IN2(keyinput115), .Q(n311) );
  XOR3X1 U329 ( .IN1(keyinput93), .IN2(N53), .IN3(n313), .Q(N737) );
  NAND2X0 U330 ( .IN1(n310), .IN2(n272), .QN(n313) );
  XOR3X1 U331 ( .IN1(keyinput92), .IN2(N49), .IN3(n314), .Q(N736) );
  NAND2X0 U332 ( .IN1(n310), .IN2(n268), .QN(n314) );
  XOR2X1 U333 ( .IN1(n315), .IN2(keyinput81), .Q(n310) );
  NAND4X0 U334 ( .IN1(n235), .IN2(n316), .IN3(n250), .IN4(n317), .QN(n315) );
  NOR2X0 U335 ( .IN1(n318), .IN2(n319), .QN(n317) );
  XOR2X1 U336 ( .IN1(keyinput58), .IN2(n253), .Q(n319) );
  XOR2X1 U337 ( .IN1(keyinput57), .IN2(n294), .Q(n318) );
  XNOR3X1 U338 ( .IN1(keyinput114), .IN2(N45), .IN3(n320), .Q(N735) );
  NAND2X0 U339 ( .IN1(n321), .IN2(n242), .QN(n320) );
  XOR3X1 U340 ( .IN1(keyinput91), .IN2(N41), .IN3(n322), .Q(N734) );
  NAND2X0 U341 ( .IN1(n321), .IN2(n246), .QN(n322) );
  XOR3X1 U342 ( .IN1(N37), .IN2(n323), .IN3(n324), .Q(N733) );
  NAND2X0 U343 ( .IN1(n321), .IN2(n272), .QN(n324) );
  XOR2X1 U344 ( .IN1(keyinput90), .IN2(keyinput113), .Q(n323) );
  XNOR3X1 U345 ( .IN1(n325), .IN2(N33), .IN3(n326), .Q(N732) );
  NAND2X0 U346 ( .IN1(n321), .IN2(n268), .QN(n326) );
  AND4X1 U347 ( .IN1(n231), .IN2(n253), .IN3(n316), .IN4(n327), .Q(n321) );
  NOR2X0 U348 ( .IN1(n298), .IN2(n328), .QN(n327) );
  XOR2X1 U349 ( .IN1(keyinput56), .IN2(n294), .Q(n328) );
  XOR2X1 U350 ( .IN1(keyinput89), .IN2(keyinput112), .Q(n325) );
  XOR3X1 U351 ( .IN1(keyinput111), .IN2(N29), .IN3(n329), .Q(N731) );
  OR2X1 U352 ( .IN1(n259), .IN2(n330), .Q(n329) );
  XOR2X1 U353 ( .IN1(N25), .IN2(n331), .Q(N730) );
  NOR2X0 U354 ( .IN1(n332), .IN2(n330), .QN(n331) );
  XOR2X1 U355 ( .IN1(N21), .IN2(n333), .Q(N729) );
  NOR2X0 U356 ( .IN1(n334), .IN2(n330), .QN(n333) );
  XOR2X1 U357 ( .IN1(N17), .IN2(n335), .Q(N728) );
  NOR2X0 U358 ( .IN1(n336), .IN2(n330), .QN(n335) );
  XOR2X1 U359 ( .IN1(n337), .IN2(keyinput80), .Q(n330) );
  NAND4X0 U360 ( .IN1(n228), .IN2(n316), .IN3(n250), .IN4(n338), .QN(n337) );
  NOR2X0 U361 ( .IN1(n294), .IN2(n339), .QN(n338) );
  XOR2X1 U362 ( .IN1(keyinput55), .IN2(n298), .Q(n339) );
  INVX0 U363 ( .INP(n235), .ZN(n298) );
  XOR3X1 U364 ( .IN1(N13), .IN2(n340), .IN3(n341), .Q(N727) );
  NAND2X0 U365 ( .IN1(n342), .IN2(n242), .QN(n341) );
  XOR2X1 U366 ( .IN1(keyinput88), .IN2(keyinput110), .Q(n340) );
  XOR3X1 U367 ( .IN1(N9), .IN2(n343), .IN3(n344), .Q(N726) );
  NAND2X0 U368 ( .IN1(n342), .IN2(n246), .QN(n344) );
  XOR2X1 U369 ( .IN1(keyinput87), .IN2(keyinput109), .Q(n343) );
  XOR3X1 U370 ( .IN1(n345), .IN2(n346), .IN3(n347), .Q(N725) );
  NAND2X0 U371 ( .IN1(n342), .IN2(n272), .QN(n347) );
  INVX0 U372 ( .INP(n348), .ZN(n342) );
  XOR2X1 U373 ( .IN1(keyinput86), .IN2(keyinput108), .Q(n345) );
  XOR3X1 U374 ( .IN1(keyinput107), .IN2(N1), .IN3(n349), .Q(N724) );
  NOR2X0 U375 ( .IN1(n336), .IN2(n348), .QN(n349) );
  NAND4X0 U376 ( .IN1(n316), .IN2(n253), .IN3(n350), .IN4(n351), .QN(n348) );
  NOR2X0 U377 ( .IN1(n352), .IN2(n294), .QN(n351) );
  INVX0 U378 ( .INP(n240), .ZN(n294) );
  XOR3X1 U379 ( .IN1(keyinput42), .IN2(keyinput38), .IN3(n353), .Q(n240) );
  XOR3X1 U380 ( .IN1(n354), .IN2(keyinput22), .IN3(n355), .Q(n353) );
  XOR3X1 U381 ( .IN1(n356), .IN2(n357), .IN3(n358), .Q(n355) );
  XOR3X1 U382 ( .IN1(n359), .IN2(n360), .IN3(n361), .Q(n358) );
  XOR2X1 U383 ( .IN1(N25), .IN2(N113), .Q(n360) );
  XOR2X1 U384 ( .IN1(n362), .IN2(n363), .Q(n357) );
  NAND2X0 U385 ( .IN1(N133), .IN2(N137), .QN(n363) );
  INVX0 U386 ( .INP(N21), .ZN(n362) );
  XOR3X1 U387 ( .IN1(N65), .IN2(N5), .IN3(n364), .Q(n356) );
  XOR2X1 U388 ( .IN1(N9), .IN2(N81), .Q(n364) );
  XOR3X1 U389 ( .IN1(keyinput21), .IN2(keyinput13), .IN3(N97), .Q(n354) );
  XOR2X1 U390 ( .IN1(n235), .IN2(keyinput53), .Q(n352) );
  XOR3X1 U391 ( .IN1(keyinput24), .IN2(keyinput14), .IN3(n365), .Q(n235) );
  XOR3X1 U392 ( .IN1(n366), .IN2(n367), .IN3(n368), .Q(n365) );
  XOR3X1 U393 ( .IN1(n369), .IN2(n370), .IN3(n371), .Q(n368) );
  XOR3X1 U394 ( .IN1(N101), .IN2(n372), .IN3(n373), .Q(n371) );
  XOR2X1 U395 ( .IN1(N37), .IN2(N117), .Q(n372) );
  XOR3X1 U396 ( .IN1(N69), .IN2(N57), .IN3(n374), .Q(n369) );
  XOR2X1 U397 ( .IN1(keyinput23), .IN2(N85), .Q(n374) );
  XOR3X1 U398 ( .IN1(keyinput33), .IN2(N53), .IN3(n375), .Q(n367) );
  XOR2X1 U399 ( .IN1(keyinput43), .IN2(keyinput39), .Q(n375) );
  XOR2X1 U400 ( .IN1(n376), .IN2(n377), .Q(n366) );
  NAND2X0 U401 ( .IN1(N134), .IN2(N137), .QN(n377) );
  XOR2X1 U402 ( .IN1(keyinput54), .IN2(n231), .Q(n350) );
  INVX0 U403 ( .INP(n250), .ZN(n231) );
  XOR3X1 U404 ( .IN1(n378), .IN2(keyinput45), .IN3(n379), .Q(n250) );
  XOR3X1 U405 ( .IN1(n380), .IN2(n381), .IN3(n382), .Q(n379) );
  XNOR2X1 U406 ( .IN1(n370), .IN2(n383), .Q(n382) );
  XNOR3X1 U407 ( .IN1(N61), .IN2(N49), .IN3(n384), .Q(n370) );
  XNOR3X1 U408 ( .IN1(keyinput4), .IN2(keyinput3), .IN3(keyinput27), .Q(n384)
         );
  INVX0 U409 ( .INP(n361), .ZN(n381) );
  XOR3X1 U410 ( .IN1(keyinput25), .IN2(keyinput0), .IN3(n385), .Q(n361) );
  XNOR2X1 U411 ( .IN1(N17), .IN2(N29), .Q(n385) );
  XOR3X1 U412 ( .IN1(keyinput32), .IN2(keyinput15), .IN3(n386), .Q(n378) );
  XNOR2X1 U413 ( .IN1(N93), .IN2(n387), .Q(n386) );
  NAND2X0 U414 ( .IN1(N136), .IN2(N137), .QN(n387) );
  INVX0 U415 ( .INP(n228), .ZN(n253) );
  XOR3X1 U416 ( .IN1(n388), .IN2(n389), .IN3(n390), .Q(n228) );
  XOR2X1 U417 ( .IN1(n373), .IN2(n359), .Q(n390) );
  XOR2X1 U418 ( .IN1(N1), .IN2(N13), .Q(n359) );
  XOR3X1 U419 ( .IN1(N45), .IN2(N33), .IN3(n391), .Q(n373) );
  XNOR3X1 U420 ( .IN1(keyinput26), .IN2(keyinput2), .IN3(keyinput1), .Q(n391)
         );
  XOR3X1 U421 ( .IN1(keyinput44), .IN2(keyinput31), .IN3(n392), .Q(n389) );
  XNOR2X1 U422 ( .IN1(N89), .IN2(n393), .Q(n392) );
  NAND2X0 U423 ( .IN1(N137), .IN2(N135), .QN(n393) );
  XOR2X1 U424 ( .IN1(n394), .IN2(n395), .Q(n388) );
  XNOR2X1 U425 ( .IN1(n396), .IN2(keyinput78), .Q(n316) );
  NAND4X0 U426 ( .IN1(n397), .IN2(n398), .IN3(n399), .IN4(n400), .QN(n396) );
  XNOR2X1 U427 ( .IN1(n401), .IN2(keyinput75), .Q(n400) );
  NAND3X0 U428 ( .IN1(n332), .IN2(n259), .IN3(n334), .QN(n401) );
  XOR2X1 U429 ( .IN1(n402), .IN2(keyinput72), .Q(n399) );
  NAND4X0 U430 ( .IN1(n242), .IN2(n403), .IN3(n404), .IN4(n405), .QN(n402) );
  XOR2X1 U431 ( .IN1(keyinput47), .IN2(n272), .Q(n405) );
  XOR2X1 U432 ( .IN1(keyinput48), .IN2(n246), .Q(n404) );
  XOR2X1 U433 ( .IN1(keyinput46), .IN2(n268), .Q(n403) );
  XOR2X1 U434 ( .IN1(n406), .IN2(keyinput73), .Q(n398) );
  NAND4X0 U435 ( .IN1(n407), .IN2(n408), .IN3(n246), .IN4(n259), .QN(n406) );
  XOR2X1 U436 ( .IN1(keyinput50), .IN2(n272), .Q(n408) );
  INVX0 U437 ( .INP(n334), .ZN(n272) );
  XOR2X1 U438 ( .IN1(keyinput49), .IN2(n268), .Q(n407) );
  XOR2X1 U439 ( .IN1(n409), .IN2(keyinput74), .Q(n397) );
  NAND3X0 U440 ( .IN1(n410), .IN2(n411), .IN3(n243), .QN(n409) );
  NOR2X0 U441 ( .IN1(n268), .IN2(n334), .QN(n243) );
  XOR3X1 U442 ( .IN1(n412), .IN2(n413), .IN3(n414), .Q(n334) );
  XOR3X1 U443 ( .IN1(n415), .IN2(n416), .IN3(n417), .Q(n414) );
  XNOR2X1 U444 ( .IN1(n383), .IN2(n394), .Q(n417) );
  XNOR3X1 U445 ( .IN1(N121), .IN2(N105), .IN3(n418), .Q(n394) );
  XOR2X1 U446 ( .IN1(N37), .IN2(n346), .Q(n418) );
  INVX0 U447 ( .INP(N5), .ZN(n346) );
  XOR3X1 U448 ( .IN1(N53), .IN2(N21), .IN3(N125), .Q(n383) );
  XOR2X1 U449 ( .IN1(keyinput18), .IN2(keyinput17), .Q(n413) );
  XOR3X1 U450 ( .IN1(keyinput35), .IN2(keyinput10), .IN3(n419), .Q(n412) );
  XOR2X1 U451 ( .IN1(n247), .IN2(n420), .Q(n419) );
  NAND2X0 U452 ( .IN1(N130), .IN2(N137), .QN(n420) );
  INVX0 U453 ( .INP(N109), .ZN(n247) );
  INVX0 U454 ( .INP(n336), .ZN(n268) );
  XOR2X1 U455 ( .IN1(keyinput51), .IN2(n246), .Q(n411) );
  INVX0 U456 ( .INP(n332), .ZN(n246) );
  XOR3X1 U457 ( .IN1(keyinput11), .IN2(N105), .IN3(n421), .Q(n332) );
  XOR3X1 U458 ( .IN1(n422), .IN2(n415), .IN3(n423), .Q(n421) );
  XNOR3X1 U459 ( .IN1(n395), .IN2(n424), .IN3(n380), .Q(n423) );
  XNOR3X1 U460 ( .IN1(N25), .IN2(N109), .IN3(n425), .Q(n380) );
  XNOR2X1 U461 ( .IN1(N57), .IN2(N77), .Q(n425) );
  XOR3X1 U462 ( .IN1(N9), .IN2(n275), .IN3(n376), .Q(n395) );
  INVX0 U463 ( .INP(N41), .ZN(n376) );
  INVX0 U464 ( .INP(N73), .ZN(n275) );
  XOR3X1 U465 ( .IN1(keyinput7), .IN2(n256), .IN3(n254), .Q(n415) );
  INVX0 U466 ( .INP(N101), .ZN(n254) );
  INVX0 U467 ( .INP(N97), .ZN(n256) );
  XNOR3X1 U468 ( .IN1(keyinput29), .IN2(keyinput19), .IN3(n426), .Q(n422) );
  NAND2X0 U469 ( .IN1(N131), .IN2(N137), .QN(n426) );
  XOR2X1 U470 ( .IN1(keyinput52), .IN2(n259), .Q(n410) );
  INVX0 U471 ( .INP(n242), .ZN(n259) );
  XOR3X1 U472 ( .IN1(n427), .IN2(n428), .IN3(n429), .Q(n242) );
  XOR3X1 U473 ( .IN1(n430), .IN2(n431), .IN3(n432), .Q(n429) );
  XOR2X1 U474 ( .IN1(n433), .IN2(n416), .Q(n432) );
  XOR3X1 U475 ( .IN1(keyinput8), .IN2(n233), .IN3(n238), .Q(n416) );
  INVX0 U476 ( .INP(N113), .ZN(n238) );
  INVX0 U477 ( .INP(N117), .ZN(n233) );
  XOR3X1 U478 ( .IN1(N13), .IN2(N125), .IN3(n434), .Q(n431) );
  XOR2X1 U479 ( .IN1(N45), .IN2(N29), .Q(n434) );
  XNOR2X1 U480 ( .IN1(N121), .IN2(n435), .Q(n430) );
  NAND2X0 U481 ( .IN1(N132), .IN2(N137), .QN(n435) );
  XOR3X1 U482 ( .IN1(keyinput30), .IN2(keyinput20), .IN3(n436), .Q(n428) );
  XOR2X1 U483 ( .IN1(keyinput41), .IN2(keyinput37), .Q(n436) );
  XOR2X1 U484 ( .IN1(keyinput12), .IN2(N61), .Q(n427) );
  XOR3X1 U485 ( .IN1(n437), .IN2(n438), .IN3(n439), .Q(n336) );
  XOR3X1 U486 ( .IN1(n440), .IN2(n441), .IN3(n442), .Q(n439) );
  XOR2X1 U487 ( .IN1(n433), .IN2(n424), .Q(n442) );
  XNOR2X1 U488 ( .IN1(N65), .IN2(n278), .Q(n424) );
  INVX0 U489 ( .INP(N69), .ZN(n278) );
  XOR3X1 U490 ( .IN1(N81), .IN2(n443), .IN3(n444), .Q(n433) );
  XOR3X1 U491 ( .IN1(keyinput6), .IN2(keyinput5), .IN3(n445), .Q(n444) );
  XNOR2X1 U492 ( .IN1(N93), .IN2(keyinput28), .Q(n445) );
  XOR2X1 U493 ( .IN1(N89), .IN2(N85), .Q(n443) );
  XOR3X1 U494 ( .IN1(N73), .IN2(N17), .IN3(n446), .Q(n441) );
  XOR2X1 U495 ( .IN1(keyinput16), .IN2(N77), .Q(n446) );
  XOR2X1 U496 ( .IN1(n447), .IN2(n448), .Q(n440) );
  NAND2X0 U497 ( .IN1(N129), .IN2(N137), .QN(n448) );
  INVX0 U498 ( .INP(N1), .ZN(n447) );
  XOR3X1 U499 ( .IN1(keyinput36), .IN2(keyinput34), .IN3(n449), .Q(n438) );
  XOR2X1 U500 ( .IN1(keyinput9), .IN2(keyinput40), .Q(n449) );
  XOR2X1 U501 ( .IN1(N49), .IN2(N33), .Q(n437) );
endmodule

