
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47,
         N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92,
         N95, N99, N102, N105, N108, N112, N115, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508;

  XNOR2X1 U256 ( .IN1(n254), .IN2(keyinput127), .Q(N432) );
  NAND3X0 U257 ( .IN1(n255), .IN2(n256), .IN3(n257), .QN(n254) );
  XOR2X1 U258 ( .IN1(n258), .IN2(keyinput124), .Q(n257) );
  NAND4X0 U259 ( .IN1(n259), .IN2(n260), .IN3(n261), .IN4(n262), .QN(n258) );
  XOR2X1 U260 ( .IN1(n263), .IN2(keyinput119), .Q(n259) );
  XNOR2X1 U261 ( .IN1(n264), .IN2(keyinput126), .Q(N431) );
  NAND4X0 U262 ( .IN1(n265), .IN2(n255), .IN3(n261), .IN4(n266), .QN(n264) );
  XOR2X1 U263 ( .IN1(n267), .IN2(keyinput122), .Q(n255) );
  NAND3X0 U264 ( .IN1(n268), .IN2(n262), .IN3(n269), .QN(n267) );
  XNOR2X1 U265 ( .IN1(keyinput117), .IN2(n270), .Q(n268) );
  XOR2X1 U266 ( .IN1(n271), .IN2(keyinput123), .Q(n265) );
  NAND3X0 U267 ( .IN1(n272), .IN2(n262), .IN3(n273), .QN(n271) );
  XNOR2X1 U268 ( .IN1(keyinput118), .IN2(n260), .Q(n273) );
  XOR2X1 U269 ( .IN1(n274), .IN2(keyinput125), .Q(N430) );
  NAND2X0 U270 ( .IN1(n256), .IN2(n269), .QN(n274) );
  AND2X1 U271 ( .IN1(n275), .IN2(n266), .Q(n256) );
  XOR2X1 U272 ( .IN1(keyinput121), .IN2(n276), .Q(n275) );
  NOR2X0 U273 ( .IN1(n277), .IN2(n278), .QN(n276) );
  XNOR2X1 U274 ( .IN1(keyinput116), .IN2(n262), .Q(n278) );
  INVX0 U275 ( .INP(n261), .ZN(n277) );
  XOR2X1 U276 ( .IN1(n279), .IN2(keyinput80), .Q(N329) );
  XOR2X1 U277 ( .IN1(keyinput120), .IN2(n280), .Q(N421) );
  NOR2X0 U278 ( .IN1(n281), .IN2(n282), .QN(n280) );
  XOR2X1 U279 ( .IN1(n283), .IN2(keyinput109), .Q(n282) );
  NAND4X0 U280 ( .IN1(N4), .IN2(n284), .IN3(n285), .IN4(n286), .QN(n283) );
  NAND2X0 U281 ( .IN1(N8), .IN2(n287), .QN(n286) );
  XOR2X1 U282 ( .IN1(keyinput101), .IN2(n288), .Q(n285) );
  NOR2X0 U283 ( .IN1(n289), .IN2(n290), .QN(n288) );
  XOR2X1 U284 ( .IN1(keyinput44), .IN2(n291), .Q(n284) );
  AND2X1 U285 ( .IN1(n292), .IN2(N1), .Q(n291) );
  XOR2X1 U286 ( .IN1(n293), .IN2(keyinput115), .Q(n281) );
  NAND4X0 U287 ( .IN1(n270), .IN2(n260), .IN3(n269), .IN4(n294), .QN(n293) );
  AND4X1 U288 ( .IN1(n262), .IN2(n263), .IN3(n295), .IN4(n266), .Q(n294) );
  XNOR2X1 U289 ( .IN1(n296), .IN2(keyinput110), .Q(n266) );
  NAND4X0 U290 ( .IN1(n297), .IN2(N17), .IN3(n298), .IN4(n299), .QN(n296) );
  NAND2X0 U291 ( .IN1(N11), .IN2(n292), .QN(n299) );
  XOR2X1 U292 ( .IN1(keyinput102), .IN2(n300), .Q(n298) );
  NOR2X0 U293 ( .IN1(n289), .IN2(n301), .QN(n300) );
  XOR2X1 U294 ( .IN1(n302), .IN2(keyinput84), .Q(n297) );
  NAND2X0 U295 ( .IN1(N21), .IN2(n287), .QN(n302) );
  OAI221X1 U296 ( .IN1(n289), .IN2(n303), .IN3(n304), .IN4(n305), .IN5(n306), 
        .QN(n295) );
  NOR2X0 U297 ( .IN1(n307), .IN2(n308), .QN(n306) );
  XOR2X1 U298 ( .IN1(keyinput53), .IN2(n309), .Q(n308) );
  AND2X1 U299 ( .IN1(n292), .IN2(N102), .Q(n309) );
  NAND4X0 U300 ( .IN1(n310), .IN2(n311), .IN3(N95), .IN4(n312), .QN(n263) );
  XOR2X1 U301 ( .IN1(keyinput92), .IN2(n313), .Q(n312) );
  AND2X1 U302 ( .IN1(n287), .IN2(N99), .Q(n313) );
  XOR2X1 U303 ( .IN1(n314), .IN2(keyinput108), .Q(n311) );
  NAND2X0 U304 ( .IN1(N105), .IN2(n315), .QN(n314) );
  XOR2X1 U305 ( .IN1(n316), .IN2(keyinput52), .Q(n310) );
  NAND2X0 U306 ( .IN1(N89), .IN2(n292), .QN(n316) );
  NAND4X0 U307 ( .IN1(n317), .IN2(n318), .IN3(N43), .IN4(n319), .QN(n262) );
  XOR2X1 U308 ( .IN1(keyinput87), .IN2(n320), .Q(n319) );
  NOR2X0 U309 ( .IN1(n304), .IN2(n321), .QN(n320) );
  XOR2X1 U310 ( .IN1(n322), .IN2(keyinput104), .Q(n318) );
  NAND2X0 U311 ( .IN1(N53), .IN2(n315), .QN(n322) );
  XOR2X1 U312 ( .IN1(n323), .IN2(keyinput48), .Q(n317) );
  NAND2X0 U313 ( .IN1(N37), .IN2(n292), .QN(n323) );
  AND2X1 U314 ( .IN1(n261), .IN2(n272), .Q(n269) );
  XNOR2X1 U315 ( .IN1(keyinput112), .IN2(n324), .Q(n272) );
  NAND4X0 U316 ( .IN1(n325), .IN2(N56), .IN3(n326), .IN4(n327), .QN(n324) );
  XOR2X1 U317 ( .IN1(keyinput49), .IN2(n328), .Q(n327) );
  AND2X1 U318 ( .IN1(n292), .IN2(N50), .Q(n328) );
  XOR2X1 U319 ( .IN1(keyinput89), .IN2(n329), .Q(n326) );
  AND2X1 U320 ( .IN1(n287), .IN2(N60), .Q(n329) );
  XOR2X1 U321 ( .IN1(n330), .IN2(keyinput105), .Q(n325) );
  NAND2X0 U322 ( .IN1(N66), .IN2(n315), .QN(n330) );
  XOR2X1 U323 ( .IN1(n331), .IN2(keyinput111), .Q(n261) );
  NAND4X0 U324 ( .IN1(n332), .IN2(N30), .IN3(n333), .IN4(n334), .QN(n331) );
  NAND2X0 U325 ( .IN1(N34), .IN2(n287), .QN(n334) );
  XOR2X1 U326 ( .IN1(keyinput103), .IN2(n335), .Q(n333) );
  AND2X1 U327 ( .IN1(n315), .IN2(N40), .Q(n335) );
  XOR2X1 U328 ( .IN1(n336), .IN2(keyinput46), .Q(n332) );
  NAND2X0 U329 ( .IN1(N24), .IN2(n292), .QN(n336) );
  XOR2X1 U330 ( .IN1(n337), .IN2(keyinput114), .Q(n260) );
  NAND4X0 U331 ( .IN1(N82), .IN2(n338), .IN3(n339), .IN4(n340), .QN(n337) );
  NAND2X0 U332 ( .IN1(N86), .IN2(n287), .QN(n340) );
  XOR2X1 U333 ( .IN1(keyinput107), .IN2(n341), .Q(n339) );
  NOR2X0 U334 ( .IN1(n289), .IN2(n342), .QN(n341) );
  INVX0 U335 ( .INP(n315), .ZN(n289) );
  XOR2X1 U336 ( .IN1(keyinput51), .IN2(n343), .Q(n338) );
  AND2X1 U337 ( .IN1(n292), .IN2(N76), .Q(n343) );
  XNOR2X1 U338 ( .IN1(keyinput113), .IN2(n344), .Q(n270) );
  NOR3X0 U339 ( .IN1(n345), .IN2(n346), .IN3(n347), .QN(n344) );
  XOR2X1 U340 ( .IN1(keyinput106), .IN2(n348), .Q(n347) );
  AND2X1 U341 ( .IN1(n315), .IN2(N79), .Q(n348) );
  XOR2X1 U342 ( .IN1(N370), .IN2(keyinput100), .Q(n315) );
  NAND4X0 U343 ( .IN1(n349), .IN2(n350), .IN3(n351), .IN4(n352), .QN(N370) );
  NOR4X0 U344 ( .IN1(n353), .IN2(n354), .IN3(n355), .IN4(n356), .QN(n352) );
  XOR2X1 U345 ( .IN1(n357), .IN2(keyinput97), .Q(n356) );
  NAND2X0 U346 ( .IN1(n358), .IN2(n359), .QN(n357) );
  XOR3X1 U347 ( .IN1(keyinput74), .IN2(keyinput67), .IN3(n360), .Q(n359) );
  NOR2X0 U348 ( .IN1(n361), .IN2(n362), .QN(n360) );
  XOR2X1 U349 ( .IN1(keyinput30), .IN2(n363), .Q(n362) );
  NOR2X0 U350 ( .IN1(N79), .IN2(n364), .QN(n363) );
  INVX0 U351 ( .INP(n365), .ZN(n361) );
  XOR3X1 U352 ( .IN1(keyinput85), .IN2(n366), .IN3(n367), .Q(n358) );
  XOR2X1 U353 ( .IN1(n368), .IN2(keyinput96), .Q(n355) );
  NAND2X0 U354 ( .IN1(n369), .IN2(n370), .QN(n368) );
  XOR2X1 U355 ( .IN1(keyinput65), .IN2(n371), .Q(n370) );
  NOR2X0 U356 ( .IN1(n372), .IN2(n373), .QN(n371) );
  XOR2X1 U357 ( .IN1(n374), .IN2(keyinput26), .Q(n373) );
  NAND2X0 U358 ( .IN1(N43), .IN2(n375), .QN(n374) );
  INVX0 U359 ( .INP(N53), .ZN(n375) );
  XOR2X1 U360 ( .IN1(n376), .IN2(n377), .Q(n369) );
  XOR2X1 U361 ( .IN1(n378), .IN2(keyinput94), .Q(n354) );
  NAND2X0 U362 ( .IN1(n379), .IN2(n380), .QN(n378) );
  XOR3X1 U363 ( .IN1(keyinput82), .IN2(n381), .IN3(n367), .Q(n380) );
  XOR2X1 U364 ( .IN1(n382), .IN2(keyinput63), .Q(n379) );
  NAND3X0 U365 ( .IN1(n383), .IN2(n301), .IN3(n384), .QN(n382) );
  XOR2X1 U366 ( .IN1(keyinput3), .IN2(N17), .Q(n384) );
  INVX0 U367 ( .INP(N27), .ZN(n301) );
  XOR2X1 U368 ( .IN1(n385), .IN2(keyinput99), .Q(n353) );
  NAND2X0 U369 ( .IN1(n386), .IN2(n387), .QN(n385) );
  XOR3X1 U370 ( .IN1(keyinput77), .IN2(keyinput70), .IN3(n388), .Q(n387) );
  NOR2X0 U371 ( .IN1(n389), .IN2(n390), .QN(n388) );
  XOR2X1 U372 ( .IN1(n391), .IN2(keyinput36), .Q(n390) );
  NAND2X0 U373 ( .IN1(n392), .IN2(n303), .QN(n391) );
  INVX0 U374 ( .INP(N115), .ZN(n303) );
  XOR3X1 U375 ( .IN1(keyinput90), .IN2(n393), .IN3(n367), .Q(n386) );
  NOR2X0 U376 ( .IN1(n394), .IN2(n395), .QN(n351) );
  XOR2X1 U377 ( .IN1(keyinput98), .IN2(n396), .Q(n395) );
  NOR2X0 U378 ( .IN1(n397), .IN2(n398), .QN(n396) );
  XOR3X1 U379 ( .IN1(keyinput88), .IN2(n399), .IN3(n377), .Q(n398) );
  XOR3X1 U380 ( .IN1(keyinput76), .IN2(keyinput69), .IN3(n400), .Q(n397) );
  NOR2X0 U381 ( .IN1(n401), .IN2(n402), .QN(n400) );
  XOR2X1 U382 ( .IN1(keyinput34), .IN2(n403), .Q(n402) );
  NOR2X0 U383 ( .IN1(N105), .IN2(n404), .QN(n403) );
  INVX0 U384 ( .INP(n405), .ZN(n401) );
  XOR2X1 U385 ( .IN1(keyinput93), .IN2(n406), .Q(n394) );
  NOR2X0 U386 ( .IN1(n407), .IN2(n408), .QN(n406) );
  XOR3X1 U387 ( .IN1(keyinput72), .IN2(keyinput55), .IN3(n409), .Q(n408) );
  NOR2X0 U388 ( .IN1(n410), .IN2(n411), .QN(n409) );
  XOR2X1 U389 ( .IN1(n412), .IN2(keyinput16), .Q(n411) );
  NAND2X0 U390 ( .IN1(n413), .IN2(n290), .QN(n412) );
  INVX0 U391 ( .INP(N14), .ZN(n290) );
  XNOR2X1 U392 ( .IN1(keyinput1), .IN2(N4), .Q(n413) );
  XOR2X1 U393 ( .IN1(n414), .IN2(n415), .Q(n410) );
  XOR3X1 U394 ( .IN1(keyinput81), .IN2(n416), .IN3(n377), .Q(n407) );
  XOR2X1 U395 ( .IN1(n417), .IN2(keyinput95), .Q(n350) );
  NAND2X0 U396 ( .IN1(n418), .IN2(n419), .QN(n417) );
  XOR2X1 U397 ( .IN1(n420), .IN2(n377), .Q(n419) );
  XOR3X1 U398 ( .IN1(keyinput73), .IN2(keyinput64), .IN3(n421), .Q(n418) );
  NAND2X0 U399 ( .IN1(n422), .IN2(n423), .QN(n421) );
  XOR2X1 U400 ( .IN1(keyinput24), .IN2(n424), .Q(n422) );
  NOR2X0 U401 ( .IN1(N40), .IN2(n425), .QN(n424) );
  MUX21X1 U402 ( .IN1(n426), .IN2(n427), .S(n377), .Q(n349) );
  INVX0 U403 ( .INP(n367), .ZN(n377) );
  XOR2X1 U404 ( .IN1(n279), .IN2(keyinput78), .Q(n367) );
  OA22X1 U405 ( .IN1(n428), .IN2(n429), .IN3(n430), .IN4(n431), .Q(n427) );
  XOR2X1 U406 ( .IN1(keyinput86), .IN2(n432), .Q(n431) );
  XNOR2X1 U407 ( .IN1(keyinput83), .IN2(n433), .Q(n429) );
  OA22X1 U408 ( .IN1(n434), .IN2(n428), .IN3(n435), .IN4(n430), .Q(n426) );
  XNOR3X1 U409 ( .IN1(keyinput75), .IN2(keyinput68), .IN3(n436), .Q(n430) );
  NAND2X0 U410 ( .IN1(n437), .IN2(n438), .QN(n436) );
  XOR2X1 U411 ( .IN1(n439), .IN2(keyinput32), .Q(n437) );
  NAND2X0 U412 ( .IN1(n440), .IN2(n342), .QN(n439) );
  INVX0 U413 ( .INP(N92), .ZN(n342) );
  XNOR2X1 U414 ( .IN1(keyinput86), .IN2(n432), .Q(n435) );
  XNOR2X1 U415 ( .IN1(n441), .IN2(keyinput66), .Q(n428) );
  NAND2X0 U416 ( .IN1(n442), .IN2(n443), .QN(n441) );
  XOR2X1 U417 ( .IN1(n444), .IN2(keyinput28), .Q(n442) );
  OR2X1 U418 ( .IN1(n445), .IN2(N66), .Q(n444) );
  XOR2X1 U419 ( .IN1(n433), .IN2(keyinput83), .Q(n434) );
  XOR2X1 U420 ( .IN1(n446), .IN2(keyinput91), .Q(n346) );
  NAND2X0 U421 ( .IN1(N73), .IN2(n287), .QN(n446) );
  INVX0 U422 ( .INP(n304), .ZN(n287) );
  XOR2X1 U423 ( .IN1(n279), .IN2(keyinput79), .Q(n304) );
  XNOR2X1 U424 ( .IN1(keyinput71), .IN2(n447), .Q(n279) );
  NOR4X0 U425 ( .IN1(n448), .IN2(n449), .IN3(n381), .IN4(n376), .QN(n447) );
  XOR2X1 U426 ( .IN1(n450), .IN2(keyinput58), .Q(n376) );
  NAND2X0 U427 ( .IN1(n451), .IN2(n452), .QN(n450) );
  INVX0 U428 ( .INP(n372), .ZN(n452) );
  XOR3X1 U429 ( .IN1(keyinput41), .IN2(n453), .IN3(n414), .Q(n372) );
  XOR2X1 U430 ( .IN1(n454), .IN2(keyinput25), .Q(n451) );
  NAND2X0 U431 ( .IN1(N43), .IN2(n321), .QN(n454) );
  INVX0 U432 ( .INP(N47), .ZN(n321) );
  XOR2X1 U433 ( .IN1(n455), .IN2(keyinput56), .Q(n381) );
  NAND2X0 U434 ( .IN1(n456), .IN2(n383), .QN(n455) );
  XOR3X1 U435 ( .IN1(keyinput39), .IN2(n457), .IN3(n414), .Q(n383) );
  XOR2X1 U436 ( .IN1(keyinput22), .IN2(n458), .Q(n456) );
  NOR2X0 U437 ( .IN1(N21), .IN2(n459), .QN(n458) );
  XNOR2X1 U438 ( .IN1(keyinput3), .IN2(N17), .Q(n459) );
  NAND3X0 U439 ( .IN1(n432), .IN2(n433), .IN3(n393), .QN(n449) );
  XNOR2X1 U440 ( .IN1(n460), .IN2(keyinput62), .Q(n393) );
  NAND2X0 U441 ( .IN1(n461), .IN2(n462), .QN(n460) );
  INVX0 U442 ( .INP(n389), .ZN(n462) );
  XOR3X1 U443 ( .IN1(keyinput47), .IN2(n463), .IN3(n414), .Q(n389) );
  XOR2X1 U444 ( .IN1(n464), .IN2(keyinput35), .Q(n461) );
  NAND2X0 U445 ( .IN1(n392), .IN2(n305), .QN(n464) );
  INVX0 U446 ( .INP(N112), .ZN(n305) );
  XOR2X1 U447 ( .IN1(n307), .IN2(keyinput13), .Q(n392) );
  INVX0 U448 ( .INP(N108), .ZN(n307) );
  NAND2X0 U449 ( .IN1(n443), .IN2(n465), .QN(n433) );
  XOR2X1 U450 ( .IN1(keyinput27), .IN2(n466), .Q(n465) );
  NOR2X0 U451 ( .IN1(N60), .IN2(n445), .QN(n466) );
  XOR2X1 U452 ( .IN1(N56), .IN2(keyinput8), .Q(n445) );
  XOR3X1 U453 ( .IN1(keyinput42), .IN2(n467), .IN3(n414), .Q(n443) );
  XNOR2X1 U454 ( .IN1(n468), .IN2(keyinput60), .Q(n432) );
  NAND2X0 U455 ( .IN1(n469), .IN2(n438), .QN(n468) );
  XOR2X1 U456 ( .IN1(n470), .IN2(n414), .Q(n438) );
  XOR2X1 U457 ( .IN1(n471), .IN2(keyinput31), .Q(n469) );
  NAND2X0 U458 ( .IN1(n440), .IN2(n472), .QN(n471) );
  INVX0 U459 ( .INP(N86), .ZN(n472) );
  XNOR2X1 U460 ( .IN1(keyinput10), .IN2(N82), .Q(n440) );
  OR4X1 U461 ( .IN1(n416), .IN2(n366), .IN3(n420), .IN4(n399), .Q(n448) );
  XNOR2X1 U462 ( .IN1(n473), .IN2(keyinput61), .Q(n399) );
  NAND2X0 U463 ( .IN1(n405), .IN2(n474), .QN(n473) );
  XOR2X1 U464 ( .IN1(keyinput33), .IN2(n475), .Q(n474) );
  NOR2X0 U465 ( .IN1(N99), .IN2(n404), .QN(n475) );
  INVX0 U466 ( .INP(N95), .ZN(n404) );
  XOR3X1 U467 ( .IN1(keyinput45), .IN2(n476), .IN3(n414), .Q(n405) );
  XNOR2X1 U468 ( .IN1(n477), .IN2(keyinput57), .Q(n420) );
  NAND2X0 U469 ( .IN1(n478), .IN2(n423), .QN(n477) );
  XNOR3X1 U470 ( .IN1(keyinput40), .IN2(n479), .IN3(n414), .Q(n423) );
  XOR2X1 U471 ( .IN1(keyinput23), .IN2(n480), .Q(n478) );
  NOR2X0 U472 ( .IN1(N34), .IN2(n425), .QN(n480) );
  XNOR2X1 U473 ( .IN1(keyinput5), .IN2(N30), .Q(n425) );
  XNOR2X1 U474 ( .IN1(n481), .IN2(keyinput59), .Q(n366) );
  NAND2X0 U475 ( .IN1(n482), .IN2(n365), .QN(n481) );
  XNOR3X1 U476 ( .IN1(keyinput43), .IN2(n483), .IN3(n414), .Q(n365) );
  XOR2X1 U477 ( .IN1(n484), .IN2(keyinput29), .Q(n482) );
  OR2X1 U478 ( .IN1(n364), .IN2(N73), .Q(n484) );
  XNOR2X1 U479 ( .IN1(n485), .IN2(keyinput54), .Q(n416) );
  NAND2X0 U480 ( .IN1(n486), .IN2(n487), .QN(n485) );
  XOR2X1 U481 ( .IN1(keyinput15), .IN2(n488), .Q(n487) );
  NOR2X0 U482 ( .IN1(N8), .IN2(n489), .QN(n488) );
  XOR2X1 U483 ( .IN1(keyinput1), .IN2(N4), .Q(n489) );
  XNOR2X1 U484 ( .IN1(n415), .IN2(n414), .Q(n486) );
  XOR2X1 U485 ( .IN1(n292), .IN2(keyinput37), .Q(n414) );
  MUX21X1 U486 ( .IN1(n490), .IN2(n491), .S(keyinput50), .Q(n345) );
  OA21X1 U487 ( .IN1(n364), .IN2(n292), .IN3(n483), .Q(n491) );
  NAND3X0 U488 ( .IN1(N69), .IN2(n292), .IN3(N63), .QN(n490) );
  INVX0 U489 ( .INP(n492), .ZN(n292) );
  XOR2X1 U490 ( .IN1(keyinput38), .IN2(n492), .Q(N223) );
  NOR4X0 U491 ( .IN1(n467), .IN2(n453), .IN3(n493), .IN4(n494), .QN(n492) );
  OR4X1 U492 ( .IN1(n415), .IN2(n479), .IN3(n463), .IN4(n476), .Q(n494) );
  XNOR2X1 U493 ( .IN1(n495), .IN2(keyinput20), .Q(n476) );
  NAND2X0 U494 ( .IN1(N95), .IN2(n496), .QN(n495) );
  XOR2X1 U495 ( .IN1(keyinput11), .IN2(N89), .Q(n496) );
  XNOR2X1 U496 ( .IN1(n497), .IN2(keyinput21), .Q(n463) );
  NAND2X0 U497 ( .IN1(N108), .IN2(n498), .QN(n497) );
  XOR2X1 U498 ( .IN1(keyinput12), .IN2(N102), .Q(n498) );
  XNOR2X1 U499 ( .IN1(n499), .IN2(keyinput17), .Q(n479) );
  NAND2X0 U500 ( .IN1(N30), .IN2(n500), .QN(n499) );
  XOR2X1 U501 ( .IN1(keyinput4), .IN2(N24), .Q(n500) );
  XNOR2X1 U502 ( .IN1(n501), .IN2(keyinput14), .Q(n415) );
  NAND2X0 U503 ( .IN1(n502), .IN2(N4), .QN(n501) );
  XNOR2X1 U504 ( .IN1(N1), .IN2(keyinput0), .Q(n502) );
  NAND3X0 U505 ( .IN1(n457), .IN2(n483), .IN3(n470), .QN(n493) );
  NAND2X0 U506 ( .IN1(n503), .IN2(N82), .QN(n470) );
  XNOR2X1 U507 ( .IN1(N76), .IN2(keyinput9), .Q(n503) );
  OR2X1 U508 ( .IN1(n364), .IN2(N63), .Q(n483) );
  INVX0 U509 ( .INP(N69), .ZN(n364) );
  NAND2X0 U510 ( .IN1(n504), .IN2(N17), .QN(n457) );
  XNOR2X1 U511 ( .IN1(N11), .IN2(keyinput2), .Q(n504) );
  XNOR2X1 U512 ( .IN1(n505), .IN2(keyinput18), .Q(n453) );
  NAND2X0 U513 ( .IN1(N43), .IN2(n506), .QN(n505) );
  XOR2X1 U514 ( .IN1(keyinput6), .IN2(N37), .Q(n506) );
  XNOR2X1 U515 ( .IN1(n507), .IN2(keyinput19), .Q(n467) );
  NAND2X0 U516 ( .IN1(N56), .IN2(n508), .QN(n507) );
  XOR2X1 U517 ( .IN1(keyinput7), .IN2(N50), .Q(n508) );
endmodule

