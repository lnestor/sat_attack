`timescale 1ns / 1ps
module c1355 (G1,G10,G11,G12,G13,G1324,G1325,G1326,G1327,G1328,G1329,G1330,
  G1331,G1332,G1333,G1334,G1335,G1336,G1337,G1338,G1339,G1340,G1341,G1342,
  G1343,G1344,G1345,G1346,G1347,G1348,G1349,G1350,G1351,G1352,G1353,G1354,
  G1355,G14,G15,G16,G17,G18,G19,G2,G20,G21,G22,G23,G24,G25,G26,G27,G28,G29,G3,
                  G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,G4,G40,G41,G5,G6,G7,G8,G9,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:66] KeyNOTWire_0;
input G1,G2,G3,G4,G5,G6,G7,G8,G9,G10,G11,G12,G13,G14,G15,G16,G17,G18,G19,G20,
  G21,G22,G23,G24,G25,G26,G27,G28,G29,G30,G31,G32,G33,G34,G35,G36,G37,G38,G39,
  G40,G41;
output G1324,G1325,G1326,G1327,G1328,G1329,G1330,G1331,G1332,G1333,G1334,G1335,
  G1336,G1337,G1338,G1339,G1340,G1341,G1342,G1343,G1344,G1345,G1346,G1347,
  G1348,G1349,G1350,G1351,G1352,G1353,G1354,G1355;

  wire G242,G245,G248,G251,G254,G257,G260,G263,G266,G269,G272,G275,G278,G281,
    G284,G287,G290,G293,G296,G299,G302,G305,G308,G311,G314,G317,G320,G323,G326,
    G329,G332,G335,G338,G341,G344,G347,G350,G353,G356,G359,G362,G363,G364,G365,
    G366,G367,G368,G369,G370,G371,G372,G373,G374,G375,G376,G377,G378,G379,G380,
    G381,G382,G383,G384,G385,G386,G387,G388,G389,G390,G391,G392,G393,G394,G395,
    G396,G397,G398,G399,G400,G401,G402,G403,G404,G405,G406,G407,G408,G409,G410,
    G411,G412,G413,G414,G415,G416,G417,G418,G419,G420,G421,G422,G423,G424,G425,
    G426,G429,G432,G435,G438,G441,G444,G447,G450,G453,G456,G459,G462,G465,G468,
    G471,G474,G477,G480,G483,G486,G489,G492,G495,G498,G501,G504,G507,G510,G513,
    G516,G519,G522,G525,G528,G531,G534,G537,G540,G543,G546,G549,G552,G555,G558,
    G561,G564,G567,G570,G571,G572,G573,G574,G575,G576,G577,G578,G579,G580,G581,
    G582,G583,G584,G585,G586,G587,G588,G589,G590,G591,G592,G593,G594,G595,G596,
    G597,G598,G599,G600,G601,G602,G607,G612,G617,G622,G627,G632,G637,G642,G645,
    G648,G651,G654,G657,G660,G663,G666,G669,G672,G675,G678,G681,G684,G687,G690,
    G691,G692,G693,G694,G695,G696,G697,G698,G699,G700,G701,G702,G703,G704,G705,
    G706,G709,G712,G715,G718,G721,G724,G727,G730,G733,G736,G739,G742,G745,G748,
    G751,G754,G755,G756,G757,G758,G759,G760,G761,G762,G763,G764,G765,G766,G767,
    G768,G769,G770,G773,G776,G779,G782,G785,G788,G791,G794,G797,G800,G803,G806,
    G809,G812,G815,G818,G819,G820,G821,G822,G823,G824,G825,G826,G827,G828,G829,
    G830,G831,G832,G833,G834,G847,G860,G873,G886,G899,G912,G925,G938,G939,G940,
    G941,G942,G943,G944,G945,G946,G947,G948,G949,G950,G951,G952,G953,G954,G955,
    G956,G957,G958,G959,G960,G961,G962,G963,G964,G965,G966,G967,G968,G969,G970,
    G971,G972,G973,G974,G975,G976,G977,G978,G979,G980,G981,G982,G983,G984,G985,
    G986,G991,G996,G1001,G1006,G1011,G1016,G1021,G1026,G1031,G1036,G1039,G1042,
    G1045,G1048,G1051,G1054,G1057,G1060,G1063,G1066,G1069,G1072,G1075,G1078,
    G1081,G1084,G1087,G1090,G1093,G1096,G1099,G1102,G1105,G1108,G1111,G1114,
    G1117,G1120,G1123,G1126,G1129,G1132,G1135,G1138,G1141,G1144,G1147,G1150,
    G1153,G1156,G1159,G1162,G1165,G1168,G1171,G1174,G1177,G1180,G1183,G1186,
    G1189,G1192,G1195,G1198,G1201,G1204,G1207,G1210,G1213,G1216,G1219,G1222,
    G1225,G1228,G1229,G1230,G1231,G1232,G1233,G1234,G1235,G1236,G1237,G1238,
    G1239,G1240,G1241,G1242,G1243,G1244,G1245,G1246,G1247,G1248,G1249,G1250,
    G1251,G1252,G1253,G1254,G1255,G1256,G1257,G1258,G1259,G1260,G1261,G1262,
    G1263,G1264,G1265,G1266,G1267,G1268,G1269,G1270,G1271,G1272,G1273,G1274,
    G1275,G1276,G1277,G1278,G1279,G1280,G1281,G1282,G1283,G1284,G1285,G1286,
    G1287,G1288,G1289,G1290,G1291,G1292,G1293,G1294,G1295,G1296,G1297,G1298,
    G1299,G1300,G1301,G1302,G1303,G1304,G1305,G1306,G1307,G1308,G1309,G1310,
    G1311,G1312,G1313,G1314,G1315,G1316,G1317,G1318,G1319,G1320,G1321,G1322,
    G1323;

  and AND2_0(G242,G33,G41);
  and AND2_1(G245,G34,G41);
  and AND2_2(G248,G35,G41);
  and AND2_3(G251,G36,G41);
  and AND2_4(G254,G37,G41);
  and AND2_5(G257,G38,G41);
  and AND2_6(G260,G39,G41);
  and AND2_7(G263,G40,G41);
  nand NAND2_0(G266,G1,G2);
  nand NAND2_1(G269,G3,G4);
  nand NAND2_2(G272,G5,G6);
  nand NAND2_3(G275,G7,G8);
  nand NAND2_4(G278,G9,G10);
  nand NAND2_5(G281,G11,G12);
  nand NAND2_6(G284,G13,G14);
  nand NAND2_7(G287,G15,G16);
  nand NAND2_8(G290,G17,G18);
  nand NAND2_9(G293,G19,G20);
  nand NAND2_10(G296,G21,G22);
  nand NAND2_11(G299,G23,G24);
  nand NAND2_12(G302,G25,G26);
  nand NAND2_13(G305,G27,G28);
  nand NAND2_14(G308,G29,G30);
  nand NAND2_15(G311,G31,G32);
  nand NAND2_16(G314,G1,G5);
  nand NAND2_17(G317,G9,G13);
  nand NAND2_18(G320,G2,G6);
  nand NAND2_19(G323,G10,G14);
  nand NAND2_20(G326,G3,G7);
  nand NAND2_21(G329,G11,G15);
  nand NAND2_22(G332,G4,G8);
  nand NAND2_23(G335,G12,G16);
  nand NAND2_24(G338,G17,G21);
  nand NAND2_25(G341,G25,G29);
  nand NAND2_26(G344,G18,G22);
  nand NAND2_27(G347,G26,G30);
  nand NAND2_28(G350,G19,G23);
  nand NAND2_29(G353,G27,G31);
  nand NAND2_30(G356,G20,G24);
  nand NAND2_31(G359,G28,G32);
  nand NAND2_32(G362,G1,G266);
  nand NAND2_33(G363,G2,G266);
  nand NAND2_34(G364,G3,G269);
  nand NAND2_35(G365,G4,G269);
  nand NAND2_36(G366,G5,G272);
  nand NAND2_37(G367,G6,G272);
  nand NAND2_38(G368,G7,G275);
  nand NAND2_39(G369,G8,G275);
  nand NAND2_40(G370,G9,G278);
  nand NAND2_41(G371,G10,G278);
  nand NAND2_42(G372,G11,G281);
  nand NAND2_43(G373,G12,G281);
  nand NAND2_44(G374,G13,G284);
  nand NAND2_45(G375,G14,G284);
  nand NAND2_46(G376,G15,G287);
  nand NAND2_47(G377,G16,G287);
  nand NAND2_48(G378,G17,G290);
  nand NAND2_49(G379,G18,G290);
  nand NAND2_50(G380,G19,G293);
  nand NAND2_51(G381,G20,G293);
  nand NAND2_52(G382,G21,G296);
  nand NAND2_53(G383,G22,G296);
  nand NAND2_54(G384,G23,G299);
  nand NAND2_55(G385,G24,G299);
  nand NAND2_56(G386,G25,G302);
  nand NAND2_57(G387,G26,G302);
  nand NAND2_58(G388,G27,G305);
  nand NAND2_59(G389,G28,G305);
  nand NAND2_60(G390,G29,G308);
  nand NAND2_61(G391,G30,G308);
  nand NAND2_62(G392,G31,G311);
  nand NAND2_63(G393,G32,G311);
  nand NAND2_64(G394,G1,G314);
  nand NAND2_65(G395,G5,G314);
  nand NAND2_66(G396,G9,G317);
  nand NAND2_67(G397,G13,G317);
  nand NAND2_68(G398,G2,G320);
  nand NAND2_69(G399,G6,G320);
  nand NAND2_70(G400,G10,G323);
  nand NAND2_71(G401,G14,G323);
  nand NAND2_72(G402,G3,G326);
  nand NAND2_73(G403,G7,G326);
  nand NAND2_74(G404,G11,G329);
  nand NAND2_75(G405,G15,G329);
  nand NAND2_76(G406,G4,G332);
  nand NAND2_77(G407,G8,G332);
  nand NAND2_78(G408,G12,G335);
  nand NAND2_79(G409,G16,G335);
  nand NAND2_80(G410,G17,G338);
  nand NAND2_81(G411,G21,G338);
  nand NAND2_82(G412,G25,G341);
  nand NAND2_83(G413,G29,G341);
  nand NAND2_84(G414,G18,G344);
  nand NAND2_85(G415,G22,G344);
  nand NAND2_86(G416,G26,G347);
  nand NAND2_87(G417,G30,G347);
  nand NAND2_88(G418,G19,G350);
  nand NAND2_89(G419,G23,G350);
  nand NAND2_90(G420,G27,G353);
  nand NAND2_91(G421,G31,G353);
  nand NAND2_92(G422,G20,G356);
  nand NAND2_93(G423,G24,G356);
  nand NAND2_94(G424,G28,G359);
  nand NAND2_95(G425,G32,G359);
  nand NAND2_96(KeyWire_0[0], G362,G363);
  xor KeyGate_0_0(G426, keyIn_0_0, KeyWire_0[0]);
  nand NAND2_97(KeyWire_0[1], G364,G365);
  xnor KeyGate_0_1(G429, keyIn_0_1, KeyWire_0[1]);
  nand NAND2_98(KeyWire_0[2], G366,G367);
  xnor KeyGate_0_2(G432, keyIn_0_2, KeyWire_0[2]);
  nand NAND2_99(KeyWire_0[3], G368,G369);
  xnor KeyGate_0_3(G435, keyIn_0_3, KeyWire_0[3]);
  nand NAND2_100(KeyWire_0[4], G370,G371);
  xnor KeyGate_0_4(G438, keyIn_0_4, KeyWire_0[4]);
  nand NAND2_101(KeyWire_0[5], G372,G373);
  xor KeyGate_0_5(KeyNOTWire_0[0], keyIn_0_5, KeyWire_0[5]);
  not KeyNOTGate_0_0(G441, KeyNOTWire_0[0]);
  nand NAND2_102(KeyWire_0[6], G374,G375);
  xnor KeyGate_0_6(G444, keyIn_0_6, KeyWire_0[6]);
  nand NAND2_103(KeyWire_0[7], G376,G377);
  xnor KeyGate_0_7(KeyNOTWire_0[1], keyIn_0_7, KeyWire_0[7]);
  not KeyNOTGate_0_1(G447, KeyNOTWire_0[1]);
  nand NAND2_104(KeyWire_0[8], G378,G379);
  xor KeyGate_0_8(KeyNOTWire_0[2], keyIn_0_8, KeyWire_0[8]);
  not KeyNOTGate_0_2(G450, KeyNOTWire_0[2]);
  nand NAND2_105(KeyWire_0[9], G380,G381);
  xnor KeyGate_0_9(KeyNOTWire_0[3], keyIn_0_9, KeyWire_0[9]);
  not KeyNOTGate_0_3(G453, KeyNOTWire_0[3]);
  nand NAND2_106(KeyWire_0[10], G382,G383);
  xor KeyGate_0_10(KeyNOTWire_0[4], keyIn_0_10, KeyWire_0[10]);
  not KeyNOTGate_0_4(G456, KeyNOTWire_0[4]);
  nand NAND2_107(KeyWire_0[11], G384,G385);
  xor KeyGate_0_11(KeyNOTWire_0[5], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_5(G459, KeyNOTWire_0[5]);
  nand NAND2_108(KeyWire_0[12], G386,G387);
  xor KeyGate_0_12(KeyNOTWire_0[6], keyIn_0_12, KeyWire_0[12]);
  not KeyNOTGate_0_6(G462, KeyNOTWire_0[6]);
  nand NAND2_109(KeyWire_0[13], G388,G389);
  xnor KeyGate_0_13(G465, keyIn_0_13, KeyWire_0[13]);
  nand NAND2_110(KeyWire_0[14], G390,G391);
  xnor KeyGate_0_14(G468, keyIn_0_14, KeyWire_0[14]);
  nand NAND2_111(KeyWire_0[15], G392,G393);
  xnor KeyGate_0_15(KeyNOTWire_0[7], keyIn_0_15, KeyWire_0[15]);
  not KeyNOTGate_0_7(G471, KeyNOTWire_0[7]);
  nand NAND2_112(KeyWire_0[16], G394,G395);
  xor KeyGate_0_16(KeyNOTWire_0[8], keyIn_0_16, KeyWire_0[16]);
  not KeyNOTGate_0_8(G474, KeyNOTWire_0[8]);
  nand NAND2_113(KeyWire_0[17], G396,G397);
  xnor KeyGate_0_17(KeyNOTWire_0[9], keyIn_0_17, KeyWire_0[17]);
  not KeyNOTGate_0_9(G477, KeyNOTWire_0[9]);
  nand NAND2_114(KeyWire_0[18], G398,G399);
  xor KeyGate_0_18(G480, keyIn_0_18, KeyWire_0[18]);
  nand NAND2_115(KeyWire_0[19], G400,G401);
  xor KeyGate_0_19(G483, keyIn_0_19, KeyWire_0[19]);
  nand NAND2_116(KeyWire_0[20], G402,G403);
  xnor KeyGate_0_20(G486, keyIn_0_20, KeyWire_0[20]);
  nand NAND2_117(KeyWire_0[21], G404,G405);
  xnor KeyGate_0_21(G489, keyIn_0_21, KeyWire_0[21]);
  nand NAND2_118(KeyWire_0[22], G406,G407);
  xor KeyGate_0_22(KeyNOTWire_0[10], keyIn_0_22, KeyWire_0[22]);
  not KeyNOTGate_0_10(G492, KeyNOTWire_0[10]);
  nand NAND2_119(KeyWire_0[23], G408,G409);
  xnor KeyGate_0_23(KeyNOTWire_0[11], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_11(G495, KeyNOTWire_0[11]);
  nand NAND2_120(KeyWire_0[24], G410,G411);
  xor KeyGate_0_24(G498, keyIn_0_24, KeyWire_0[24]);
  nand NAND2_121(KeyWire_0[25], G412,G413);
  xnor KeyGate_0_25(KeyNOTWire_0[12], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_12(G501, KeyNOTWire_0[12]);
  nand NAND2_122(KeyWire_0[26], G414,G415);
  xor KeyGate_0_26(KeyNOTWire_0[13], keyIn_0_26, KeyWire_0[26]);
  not KeyNOTGate_0_13(G504, KeyNOTWire_0[13]);
  nand NAND2_123(KeyWire_0[27], G416,G417);
  xor KeyGate_0_27(KeyNOTWire_0[14], keyIn_0_27, KeyWire_0[27]);
  not KeyNOTGate_0_14(G507, KeyNOTWire_0[14]);
  nand NAND2_124(KeyWire_0[28], G418,G419);
  xor KeyGate_0_28(KeyNOTWire_0[15], keyIn_0_28, KeyWire_0[28]);
  not KeyNOTGate_0_15(G510, KeyNOTWire_0[15]);
  nand NAND2_125(KeyWire_0[29], G420,G421);
  xor KeyGate_0_29(G513, keyIn_0_29, KeyWire_0[29]);
  nand NAND2_126(KeyWire_0[30], G422,G423);
  xor KeyGate_0_30(KeyNOTWire_0[16], keyIn_0_30, KeyWire_0[30]);
  not KeyNOTGate_0_16(G516, KeyNOTWire_0[16]);
  nand NAND2_127(KeyWire_0[31], G424,G425);
  xnor KeyGate_0_31(G519, keyIn_0_31, KeyWire_0[31]);
  nand NAND2_128(KeyWire_0[32], G426,G429);
  xnor KeyGate_0_32(KeyNOTWire_0[17], keyIn_0_32, KeyWire_0[32]);
  not KeyNOTGate_0_17(G522, KeyNOTWire_0[17]);
  nand NAND2_129(KeyWire_0[33], G432,G435);
  xor KeyGate_0_33(KeyNOTWire_0[18], keyIn_0_33, KeyWire_0[33]);
  not KeyNOTGate_0_18(G525, KeyNOTWire_0[18]);
  nand NAND2_130(KeyWire_0[34], G438,G441);
  xor KeyGate_0_34(KeyNOTWire_0[19], keyIn_0_34, KeyWire_0[34]);
  not KeyNOTGate_0_19(G528, KeyNOTWire_0[19]);
  nand NAND2_131(KeyWire_0[35], G444,G447);
  xnor KeyGate_0_35(G531, keyIn_0_35, KeyWire_0[35]);
  nand NAND2_132(KeyWire_0[36], G450,G453);
  xor KeyGate_0_36(G534, keyIn_0_36, KeyWire_0[36]);
  nand NAND2_133(KeyWire_0[37], G456,G459);
  xnor KeyGate_0_37(G537, keyIn_0_37, KeyWire_0[37]);
  nand NAND2_134(KeyWire_0[38], G462,G465);
  xor KeyGate_0_38(KeyNOTWire_0[20], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_20(G540, KeyNOTWire_0[20]);
  nand NAND2_135(KeyWire_0[39], G468,G471);
  xor KeyGate_0_39(KeyNOTWire_0[21], keyIn_0_39, KeyWire_0[39]);
  not KeyNOTGate_0_21(G543, KeyNOTWire_0[21]);
  nand NAND2_136(KeyWire_0[40], G474,G477);
  xor KeyGate_0_40(G546, keyIn_0_40, KeyWire_0[40]);
  nand NAND2_137(KeyWire_0[41], G480,G483);
  xor KeyGate_0_41(KeyNOTWire_0[22], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_22(G549, KeyNOTWire_0[22]);
  nand NAND2_138(KeyWire_0[42], G486,G489);
  xnor KeyGate_0_42(KeyNOTWire_0[23], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_23(G552, KeyNOTWire_0[23]);
  nand NAND2_139(KeyWire_0[43], G492,G495);
  xnor KeyGate_0_43(G555, keyIn_0_43, KeyWire_0[43]);
  nand NAND2_140(KeyWire_0[44], G498,G501);
  xor KeyGate_0_44(G558, keyIn_0_44, KeyWire_0[44]);
  nand NAND2_141(KeyWire_0[45], G504,G507);
  xor KeyGate_0_45(G561, keyIn_0_45, KeyWire_0[45]);
  nand NAND2_142(KeyWire_0[46], G510,G513);
  xnor KeyGate_0_46(KeyNOTWire_0[24], keyIn_0_46, KeyWire_0[46]);
  not KeyNOTGate_0_24(G564, KeyNOTWire_0[24]);
  nand NAND2_143(KeyWire_0[47], G516,G519);
  xor KeyGate_0_47(G567, keyIn_0_47, KeyWire_0[47]);
  nand NAND2_144(KeyWire_0[48], G426,G522);
  xor KeyGate_0_48(G570, keyIn_0_48, KeyWire_0[48]);
  nand NAND2_145(KeyWire_0[49], G429,G522);
  xnor KeyGate_0_49(KeyNOTWire_0[25], keyIn_0_49, KeyWire_0[49]);
  not KeyNOTGate_0_25(G571, KeyNOTWire_0[25]);
  nand NAND2_146(KeyWire_0[50], G432,G525);
  xnor KeyGate_0_50(G572, keyIn_0_50, KeyWire_0[50]);
  nand NAND2_147(KeyWire_0[51], G435,G525);
  xor KeyGate_0_51(G573, keyIn_0_51, KeyWire_0[51]);
  nand NAND2_148(KeyWire_0[52], G438,G528);
  xnor KeyGate_0_52(KeyNOTWire_0[26], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_26(G574, KeyNOTWire_0[26]);
  nand NAND2_149(KeyWire_0[53], G441,G528);
  xor KeyGate_0_53(KeyNOTWire_0[27], keyIn_0_53, KeyWire_0[53]);
  not KeyNOTGate_0_27(G575, KeyNOTWire_0[27]);
  nand NAND2_150(KeyWire_0[54], G444,G531);
  xor KeyGate_0_54(G576, keyIn_0_54, KeyWire_0[54]);
  nand NAND2_151(KeyWire_0[55], G447,G531);
  xor KeyGate_0_55(KeyNOTWire_0[28], keyIn_0_55, KeyWire_0[55]);
  not KeyNOTGate_0_28(G577, KeyNOTWire_0[28]);
  nand NAND2_152(KeyWire_0[56], G450,G534);
  xor KeyGate_0_56(KeyNOTWire_0[29], keyIn_0_56, KeyWire_0[56]);
  not KeyNOTGate_0_29(G578, KeyNOTWire_0[29]);
  nand NAND2_153(KeyWire_0[57], G453,G534);
  xor KeyGate_0_57(KeyNOTWire_0[30], keyIn_0_57, KeyWire_0[57]);
  not KeyNOTGate_0_30(G579, KeyNOTWire_0[30]);
  nand NAND2_154(KeyWire_0[58], G456,G537);
  xor KeyGate_0_58(KeyNOTWire_0[31], keyIn_0_58, KeyWire_0[58]);
  not KeyNOTGate_0_31(G580, KeyNOTWire_0[31]);
  nand NAND2_155(KeyWire_0[59], G459,G537);
  xor KeyGate_0_59(KeyNOTWire_0[32], keyIn_0_59, KeyWire_0[59]);
  not KeyNOTGate_0_32(G581, KeyNOTWire_0[32]);
  nand NAND2_156(KeyWire_0[60], G462,G540);
  xor KeyGate_0_60(G582, keyIn_0_60, KeyWire_0[60]);
  nand NAND2_157(KeyWire_0[61], G465,G540);
  xor KeyGate_0_61(KeyNOTWire_0[33], keyIn_0_61, KeyWire_0[61]);
  not KeyNOTGate_0_33(G583, KeyNOTWire_0[33]);
  nand NAND2_158(KeyWire_0[62], G468,G543);
  xnor KeyGate_0_62(KeyNOTWire_0[34], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_34(G584, KeyNOTWire_0[34]);
  nand NAND2_159(KeyWire_0[63], G471,G543);
  xor KeyGate_0_63(KeyNOTWire_0[35], keyIn_0_63, KeyWire_0[63]);
  not KeyNOTGate_0_35(G585, KeyNOTWire_0[35]);
  nand NAND2_160(KeyWire_0[64], G474,G546);
  xnor KeyGate_0_64(KeyNOTWire_0[36], keyIn_0_64, KeyWire_0[64]);
  not KeyNOTGate_0_36(G586, KeyNOTWire_0[36]);
  nand NAND2_161(KeyWire_0[65], G477,G546);
  xor KeyGate_0_65(G587, keyIn_0_65, KeyWire_0[65]);
  nand NAND2_162(KeyWire_0[66], G480,G549);
  xor KeyGate_0_66(KeyNOTWire_0[37], keyIn_0_66, KeyWire_0[66]);
  not KeyNOTGate_0_37(G588, KeyNOTWire_0[37]);
  nand NAND2_163(KeyWire_0[67], G483,G549);
  xnor KeyGate_0_67(KeyNOTWire_0[38], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_38(G589, KeyNOTWire_0[38]);
  nand NAND2_164(KeyWire_0[68], G486,G552);
  xor KeyGate_0_68(G590, keyIn_0_68, KeyWire_0[68]);
  nand NAND2_165(KeyWire_0[69], G489,G552);
  xnor KeyGate_0_69(G591, keyIn_0_69, KeyWire_0[69]);
  nand NAND2_166(KeyWire_0[70], G492,G555);
  xnor KeyGate_0_70(G592, keyIn_0_70, KeyWire_0[70]);
  nand NAND2_167(KeyWire_0[71], G495,G555);
  xor KeyGate_0_71(G593, keyIn_0_71, KeyWire_0[71]);
  nand NAND2_168(KeyWire_0[72], G498,G558);
  xnor KeyGate_0_72(G594, keyIn_0_72, KeyWire_0[72]);
  nand NAND2_169(KeyWire_0[73], G501,G558);
  xor KeyGate_0_73(G595, keyIn_0_73, KeyWire_0[73]);
  nand NAND2_170(KeyWire_0[74], G504,G561);
  xor KeyGate_0_74(KeyNOTWire_0[39], keyIn_0_74, KeyWire_0[74]);
  not KeyNOTGate_0_39(G596, KeyNOTWire_0[39]);
  nand NAND2_171(KeyWire_0[75], G507,G561);
  xor KeyGate_0_75(KeyNOTWire_0[40], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_40(G597, KeyNOTWire_0[40]);
  nand NAND2_172(KeyWire_0[76], G510,G564);
  xnor KeyGate_0_76(KeyNOTWire_0[41], keyIn_0_76, KeyWire_0[76]);
  not KeyNOTGate_0_41(G598, KeyNOTWire_0[41]);
  nand NAND2_173(KeyWire_0[77], G513,G564);
  xnor KeyGate_0_77(G599, keyIn_0_77, KeyWire_0[77]);
  nand NAND2_174(KeyWire_0[78], G516,G567);
  xnor KeyGate_0_78(G600, keyIn_0_78, KeyWire_0[78]);
  nand NAND2_175(KeyWire_0[79], G519,G567);
  xnor KeyGate_0_79(G601, keyIn_0_79, KeyWire_0[79]);
  nand NAND2_176(KeyWire_0[80], G570,G571);
  xnor KeyGate_0_80(KeyNOTWire_0[42], keyIn_0_80, KeyWire_0[80]);
  not KeyNOTGate_0_42(G602, KeyNOTWire_0[42]);
  nand NAND2_177(KeyWire_0[81], G572,G573);
  xnor KeyGate_0_81(G607, keyIn_0_81, KeyWire_0[81]);
  nand NAND2_178(KeyWire_0[82], G574,G575);
  xnor KeyGate_0_82(G612, keyIn_0_82, KeyWire_0[82]);
  nand NAND2_179(KeyWire_0[83], G576,G577);
  xnor KeyGate_0_83(KeyNOTWire_0[43], keyIn_0_83, KeyWire_0[83]);
  not KeyNOTGate_0_43(G617, KeyNOTWire_0[43]);
  nand NAND2_180(KeyWire_0[84], G578,G579);
  xnor KeyGate_0_84(KeyNOTWire_0[44], keyIn_0_84, KeyWire_0[84]);
  not KeyNOTGate_0_44(G622, KeyNOTWire_0[44]);
  nand NAND2_181(KeyWire_0[85], G580,G581);
  xnor KeyGate_0_85(G627, keyIn_0_85, KeyWire_0[85]);
  nand NAND2_182(KeyWire_0[86], G582,G583);
  xor KeyGate_0_86(G632, keyIn_0_86, KeyWire_0[86]);
  nand NAND2_183(KeyWire_0[87], G584,G585);
  xnor KeyGate_0_87(G637, keyIn_0_87, KeyWire_0[87]);
  nand NAND2_184(G642,G586,G587);
  nand NAND2_185(G645,G588,G589);
  nand NAND2_186(G648,G590,G591);
  nand NAND2_187(G651,G592,G593);
  nand NAND2_188(G654,G594,G595);
  nand NAND2_189(G657,G596,G597);
  nand NAND2_190(G660,G598,G599);
  nand NAND2_191(G663,G600,G601);
  nand NAND2_192(KeyWire_0[88], G602,G607);
  xnor KeyGate_0_88(G666, keyIn_0_88, KeyWire_0[88]);
  nand NAND2_193(KeyWire_0[89], G612,G617);
  xor KeyGate_0_89(G669, keyIn_0_89, KeyWire_0[89]);
  nand NAND2_194(KeyWire_0[90], G602,G612);
  xor KeyGate_0_90(G672, keyIn_0_90, KeyWire_0[90]);
  nand NAND2_195(KeyWire_0[91], G607,G617);
  xor KeyGate_0_91(KeyNOTWire_0[45], keyIn_0_91, KeyWire_0[91]);
  not KeyNOTGate_0_45(G675, KeyNOTWire_0[45]);
  nand NAND2_196(KeyWire_0[92], G622,G627);
  xnor KeyGate_0_92(KeyNOTWire_0[46], keyIn_0_92, KeyWire_0[92]);
  not KeyNOTGate_0_46(G678, KeyNOTWire_0[46]);
  nand NAND2_197(KeyWire_0[93], G632,G637);
  xnor KeyGate_0_93(KeyNOTWire_0[47], keyIn_0_93, KeyWire_0[93]);
  not KeyNOTGate_0_47(G681, KeyNOTWire_0[47]);
  nand NAND2_198(KeyWire_0[94], G622,G632);
  xnor KeyGate_0_94(KeyNOTWire_0[48], keyIn_0_94, KeyWire_0[94]);
  not KeyNOTGate_0_48(G684, KeyNOTWire_0[48]);
  nand NAND2_199(KeyWire_0[95], G627,G637);
  xnor KeyGate_0_95(KeyNOTWire_0[49], keyIn_0_95, KeyWire_0[95]);
  not KeyNOTGate_0_49(G687, KeyNOTWire_0[49]);
  nand NAND2_200(KeyWire_0[96], G602,G666);
  xnor KeyGate_0_96(G690, keyIn_0_96, KeyWire_0[96]);
  nand NAND2_201(KeyWire_0[97], G607,G666);
  xnor KeyGate_0_97(KeyNOTWire_0[50], keyIn_0_97, KeyWire_0[97]);
  not KeyNOTGate_0_50(G691, KeyNOTWire_0[50]);
  nand NAND2_202(KeyWire_0[98], G612,G669);
  xor KeyGate_0_98(G692, keyIn_0_98, KeyWire_0[98]);
  nand NAND2_203(KeyWire_0[99], G617,G669);
  xnor KeyGate_0_99(G693, keyIn_0_99, KeyWire_0[99]);
  nand NAND2_204(KeyWire_0[100], G602,G672);
  xor KeyGate_0_100(KeyNOTWire_0[51], keyIn_0_100, KeyWire_0[100]);
  not KeyNOTGate_0_51(G694, KeyNOTWire_0[51]);
  nand NAND2_205(KeyWire_0[101], G612,G672);
  xnor KeyGate_0_101(G695, keyIn_0_101, KeyWire_0[101]);
  nand NAND2_206(KeyWire_0[102], G607,G675);
  xnor KeyGate_0_102(G696, keyIn_0_102, KeyWire_0[102]);
  nand NAND2_207(KeyWire_0[103], G617,G675);
  xor KeyGate_0_103(KeyNOTWire_0[52], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_52(G697, KeyNOTWire_0[52]);
  nand NAND2_208(KeyWire_0[104], G622,G678);
  xor KeyGate_0_104(G698, keyIn_0_104, KeyWire_0[104]);
  nand NAND2_209(KeyWire_0[105], G627,G678);
  xor KeyGate_0_105(KeyNOTWire_0[53], keyIn_0_105, KeyWire_0[105]);
  not KeyNOTGate_0_53(G699, KeyNOTWire_0[53]);
  nand NAND2_210(KeyWire_0[106], G632,G681);
  xnor KeyGate_0_106(G700, keyIn_0_106, KeyWire_0[106]);
  nand NAND2_211(KeyWire_0[107], G637,G681);
  xnor KeyGate_0_107(KeyNOTWire_0[54], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_54(G701, KeyNOTWire_0[54]);
  nand NAND2_212(KeyWire_0[108], G622,G684);
  xor KeyGate_0_108(G702, keyIn_0_108, KeyWire_0[108]);
  nand NAND2_213(KeyWire_0[109], G632,G684);
  xor KeyGate_0_109(KeyNOTWire_0[55], keyIn_0_109, KeyWire_0[109]);
  not KeyNOTGate_0_55(G703, KeyNOTWire_0[55]);
  nand NAND2_214(KeyWire_0[110], G627,G687);
  xnor KeyGate_0_110(G704, keyIn_0_110, KeyWire_0[110]);
  nand NAND2_215(KeyWire_0[111], G637,G687);
  xnor KeyGate_0_111(KeyNOTWire_0[56], keyIn_0_111, KeyWire_0[111]);
  not KeyNOTGate_0_56(G705, KeyNOTWire_0[56]);
  nand NAND2_216(KeyWire_0[112], G690,G691);
  xor KeyGate_0_112(G706, keyIn_0_112, KeyWire_0[112]);
  nand NAND2_217(KeyWire_0[113], G692,G693);
  xor KeyGate_0_113(KeyNOTWire_0[57], keyIn_0_113, KeyWire_0[113]);
  not KeyNOTGate_0_57(G709, KeyNOTWire_0[57]);
  nand NAND2_218(KeyWire_0[114], G694,G695);
  xor KeyGate_0_114(KeyNOTWire_0[58], keyIn_0_114, KeyWire_0[114]);
  not KeyNOTGate_0_58(G712, KeyNOTWire_0[58]);
  nand NAND2_219(KeyWire_0[115], G696,G697);
  xnor KeyGate_0_115(KeyNOTWire_0[59], keyIn_0_115, KeyWire_0[115]);
  not KeyNOTGate_0_59(G715, KeyNOTWire_0[59]);
  nand NAND2_220(KeyWire_0[116], G698,G699);
  xor KeyGate_0_116(KeyNOTWire_0[60], keyIn_0_116, KeyWire_0[116]);
  not KeyNOTGate_0_60(G718, KeyNOTWire_0[60]);
  nand NAND2_221(KeyWire_0[117], G700,G701);
  xor KeyGate_0_117(G721, keyIn_0_117, KeyWire_0[117]);
  nand NAND2_222(KeyWire_0[118], G702,G703);
  xnor KeyGate_0_118(G724, keyIn_0_118, KeyWire_0[118]);
  nand NAND2_223(KeyWire_0[119], G704,G705);
  xor KeyGate_0_119(G727, keyIn_0_119, KeyWire_0[119]);
  nand NAND2_224(KeyWire_0[120], G242,G718);
  xnor KeyGate_0_120(G730, keyIn_0_120, KeyWire_0[120]);
  nand NAND2_225(KeyWire_0[121], G245,G721);
  xor KeyGate_0_121(KeyNOTWire_0[61], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_61(G733, KeyNOTWire_0[61]);
  nand NAND2_226(KeyWire_0[122], G248,G724);
  xnor KeyGate_0_122(KeyNOTWire_0[62], keyIn_0_122, KeyWire_0[122]);
  not KeyNOTGate_0_62(G736, KeyNOTWire_0[62]);
  nand NAND2_227(KeyWire_0[123], G251,G727);
  xnor KeyGate_0_123(KeyNOTWire_0[63], keyIn_0_123, KeyWire_0[123]);
  not KeyNOTGate_0_63(G739, KeyNOTWire_0[63]);
  nand NAND2_228(KeyWire_0[124], G254,G706);
  xnor KeyGate_0_124(KeyNOTWire_0[64], keyIn_0_124, KeyWire_0[124]);
  not KeyNOTGate_0_64(G742, KeyNOTWire_0[64]);
  nand NAND2_229(KeyWire_0[125], G257,G709);
  xnor KeyGate_0_125(KeyNOTWire_0[65], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_65(G745, KeyNOTWire_0[65]);
  nand NAND2_230(KeyWire_0[126], G260,G712);
  xor KeyGate_0_126(KeyNOTWire_0[66], keyIn_0_126, KeyWire_0[126]);
  not KeyNOTGate_0_66(G748, KeyNOTWire_0[66]);
  nand NAND2_231(KeyWire_0[127], G263,G715);
  xnor KeyGate_0_127(G751, keyIn_0_127, KeyWire_0[127]);
  nand NAND2_232(G754,G242,G730);
  nand NAND2_233(G755,G718,G730);
  nand NAND2_234(G756,G245,G733);
  nand NAND2_235(G757,G721,G733);
  nand NAND2_236(G758,G248,G736);
  nand NAND2_237(G759,G724,G736);
  nand NAND2_238(G760,G251,G739);
  nand NAND2_239(G761,G727,G739);
  nand NAND2_240(G762,G254,G742);
  nand NAND2_241(G763,G706,G742);
  nand NAND2_242(G764,G257,G745);
  nand NAND2_243(G765,G709,G745);
  nand NAND2_244(G766,G260,G748);
  nand NAND2_245(G767,G712,G748);
  nand NAND2_246(G768,G263,G751);
  nand NAND2_247(G769,G715,G751);
  nand NAND2_248(G770,G754,G755);
  nand NAND2_249(G773,G756,G757);
  nand NAND2_250(G776,G758,G759);
  nand NAND2_251(G779,G760,G761);
  nand NAND2_252(G782,G762,G763);
  nand NAND2_253(G785,G764,G765);
  nand NAND2_254(G788,G766,G767);
  nand NAND2_255(G791,G768,G769);
  nand NAND2_256(G794,G642,G770);
  nand NAND2_257(G797,G645,G773);
  nand NAND2_258(G800,G648,G776);
  nand NAND2_259(G803,G651,G779);
  nand NAND2_260(G806,G654,G782);
  nand NAND2_261(G809,G657,G785);
  nand NAND2_262(G812,G660,G788);
  nand NAND2_263(G815,G663,G791);
  nand NAND2_264(G818,G642,G794);
  nand NAND2_265(G819,G770,G794);
  nand NAND2_266(G820,G645,G797);
  nand NAND2_267(G821,G773,G797);
  nand NAND2_268(G822,G648,G800);
  nand NAND2_269(G823,G776,G800);
  nand NAND2_270(G824,G651,G803);
  nand NAND2_271(G825,G779,G803);
  nand NAND2_272(G826,G654,G806);
  nand NAND2_273(G827,G782,G806);
  nand NAND2_274(G828,G657,G809);
  nand NAND2_275(G829,G785,G809);
  nand NAND2_276(G830,G660,G812);
  nand NAND2_277(G831,G788,G812);
  nand NAND2_278(G832,G663,G815);
  nand NAND2_279(G833,G791,G815);
  nand NAND2_280(G834,G818,G819);
  nand NAND2_281(G847,G820,G821);
  nand NAND2_282(G860,G822,G823);
  nand NAND2_283(G873,G824,G825);
  nand NAND2_284(G886,G828,G829);
  nand NAND2_285(G899,G832,G833);
  nand NAND2_286(G912,G830,G831);
  nand NAND2_287(G925,G826,G827);
  not NOT_0(G938,G834);
  not NOT_1(G939,G847);
  not NOT_2(G940,G860);
  not NOT_3(G941,G834);
  not NOT_4(G942,G847);
  not NOT_5(G943,G873);
  not NOT_6(G944,G834);
  not NOT_7(G945,G860);
  not NOT_8(G946,G873);
  not NOT_9(G947,G847);
  not NOT_10(G948,G860);
  not NOT_11(G949,G873);
  not NOT_12(G950,G886);
  not NOT_13(G951,G899);
  not NOT_14(G952,G886);
  not NOT_15(G953,G912);
  not NOT_16(G954,G925);
  not NOT_17(G955,G899);
  not NOT_18(G956,G925);
  not NOT_19(G957,G912);
  not NOT_20(G958,G925);
  not NOT_21(G959,G886);
  not NOT_22(G960,G912);
  not NOT_23(G961,G925);
  not NOT_24(G962,G886);
  not NOT_25(G963,G899);
  not NOT_26(G964,G925);
  not NOT_27(G965,G912);
  not NOT_28(G966,G899);
  not NOT_29(G967,G886);
  not NOT_30(G968,G912);
  not NOT_31(G969,G899);
  not NOT_32(G970,G847);
  not NOT_33(G971,G873);
  not NOT_34(G972,G847);
  not NOT_35(G973,G860);
  not NOT_36(G974,G834);
  not NOT_37(G975,G873);
  not NOT_38(G976,G834);
  not NOT_39(G977,G860);
  and AND4_0(G978,G938,G939,G940,G873);
  and AND4_1(G979,G941,G942,G860,G943);
  and AND4_2(G980,G944,G847,G945,G946);
  and AND4_3(G981,G834,G947,G948,G949);
  and AND4_4(G982,G958,G959,G960,G899);
  and AND4_5(G983,G961,G962,G912,G963);
  and AND4_6(G984,G964,G886,G965,G966);
  and AND4_7(G985,G925,G967,G968,G969);
  or OR4_0(G986,G978,G979,G980,G981);
  or OR4_1(G991,G982,G983,G984,G985);
  and AND5_0(G996,G925,G950,G912,G951,G986);
  and AND5_1(G1001,G925,G952,G953,G899,G986);
  and AND5_2(G1006,G954,G886,G912,G955,G986);
  and AND5_3(G1011,G956,G886,G957,G899,G986);
  and AND5_4(G1016,G834,G970,G860,G971,G991);
  and AND5_5(G1021,G834,G972,G973,G873,G991);
  and AND5_6(G1026,G974,G847,G860,G975,G991);
  and AND5_7(G1031,G976,G847,G977,G873,G991);
  and AND2_8(G1036,G834,G996);
  and AND2_9(G1039,G847,G996);
  and AND2_10(G1042,G860,G996);
  and AND2_11(G1045,G873,G996);
  and AND2_12(G1048,G834,G1001);
  and AND2_13(G1051,G847,G1001);
  and AND2_14(G1054,G860,G1001);
  and AND2_15(G1057,G873,G1001);
  and AND2_16(G1060,G834,G1006);
  and AND2_17(G1063,G847,G1006);
  and AND2_18(G1066,G860,G1006);
  and AND2_19(G1069,G873,G1006);
  and AND2_20(G1072,G834,G1011);
  and AND2_21(G1075,G847,G1011);
  and AND2_22(G1078,G860,G1011);
  and AND2_23(G1081,G873,G1011);
  and AND2_24(G1084,G925,G1016);
  and AND2_25(G1087,G886,G1016);
  and AND2_26(G1090,G912,G1016);
  and AND2_27(G1093,G899,G1016);
  and AND2_28(G1096,G925,G1021);
  and AND2_29(G1099,G886,G1021);
  and AND2_30(G1102,G912,G1021);
  and AND2_31(G1105,G899,G1021);
  and AND2_32(G1108,G925,G1026);
  and AND2_33(G1111,G886,G1026);
  and AND2_34(G1114,G912,G1026);
  and AND2_35(G1117,G899,G1026);
  and AND2_36(G1120,G925,G1031);
  and AND2_37(G1123,G886,G1031);
  and AND2_38(G1126,G912,G1031);
  and AND2_39(G1129,G899,G1031);
  nand NAND2_288(G1132,G1,G1036);
  nand NAND2_289(G1135,G2,G1039);
  nand NAND2_290(G1138,G3,G1042);
  nand NAND2_291(G1141,G4,G1045);
  nand NAND2_292(G1144,G5,G1048);
  nand NAND2_293(G1147,G6,G1051);
  nand NAND2_294(G1150,G7,G1054);
  nand NAND2_295(G1153,G8,G1057);
  nand NAND2_296(G1156,G9,G1060);
  nand NAND2_297(G1159,G10,G1063);
  nand NAND2_298(G1162,G11,G1066);
  nand NAND2_299(G1165,G12,G1069);
  nand NAND2_300(G1168,G13,G1072);
  nand NAND2_301(G1171,G14,G1075);
  nand NAND2_302(G1174,G15,G1078);
  nand NAND2_303(G1177,G16,G1081);
  nand NAND2_304(G1180,G17,G1084);
  nand NAND2_305(G1183,G18,G1087);
  nand NAND2_306(G1186,G19,G1090);
  nand NAND2_307(G1189,G20,G1093);
  nand NAND2_308(G1192,G21,G1096);
  nand NAND2_309(G1195,G22,G1099);
  nand NAND2_310(G1198,G23,G1102);
  nand NAND2_311(G1201,G24,G1105);
  nand NAND2_312(G1204,G25,G1108);
  nand NAND2_313(G1207,G26,G1111);
  nand NAND2_314(G1210,G27,G1114);
  nand NAND2_315(G1213,G28,G1117);
  nand NAND2_316(G1216,G29,G1120);
  nand NAND2_317(G1219,G30,G1123);
  nand NAND2_318(G1222,G31,G1126);
  nand NAND2_319(G1225,G32,G1129);
  nand NAND2_320(G1228,G1,G1132);
  nand NAND2_321(G1229,G1036,G1132);
  nand NAND2_322(G1230,G2,G1135);
  nand NAND2_323(G1231,G1039,G1135);
  nand NAND2_324(G1232,G3,G1138);
  nand NAND2_325(G1233,G1042,G1138);
  nand NAND2_326(G1234,G4,G1141);
  nand NAND2_327(G1235,G1045,G1141);
  nand NAND2_328(G1236,G5,G1144);
  nand NAND2_329(G1237,G1048,G1144);
  nand NAND2_330(G1238,G6,G1147);
  nand NAND2_331(G1239,G1051,G1147);
  nand NAND2_332(G1240,G7,G1150);
  nand NAND2_333(G1241,G1054,G1150);
  nand NAND2_334(G1242,G8,G1153);
  nand NAND2_335(G1243,G1057,G1153);
  nand NAND2_336(G1244,G9,G1156);
  nand NAND2_337(G1245,G1060,G1156);
  nand NAND2_338(G1246,G10,G1159);
  nand NAND2_339(G1247,G1063,G1159);
  nand NAND2_340(G1248,G11,G1162);
  nand NAND2_341(G1249,G1066,G1162);
  nand NAND2_342(G1250,G12,G1165);
  nand NAND2_343(G1251,G1069,G1165);
  nand NAND2_344(G1252,G13,G1168);
  nand NAND2_345(G1253,G1072,G1168);
  nand NAND2_346(G1254,G14,G1171);
  nand NAND2_347(G1255,G1075,G1171);
  nand NAND2_348(G1256,G15,G1174);
  nand NAND2_349(G1257,G1078,G1174);
  nand NAND2_350(G1258,G16,G1177);
  nand NAND2_351(G1259,G1081,G1177);
  nand NAND2_352(G1260,G17,G1180);
  nand NAND2_353(G1261,G1084,G1180);
  nand NAND2_354(G1262,G18,G1183);
  nand NAND2_355(G1263,G1087,G1183);
  nand NAND2_356(G1264,G19,G1186);
  nand NAND2_357(G1265,G1090,G1186);
  nand NAND2_358(G1266,G20,G1189);
  nand NAND2_359(G1267,G1093,G1189);
  nand NAND2_360(G1268,G21,G1192);
  nand NAND2_361(G1269,G1096,G1192);
  nand NAND2_362(G1270,G22,G1195);
  nand NAND2_363(G1271,G1099,G1195);
  nand NAND2_364(G1272,G23,G1198);
  nand NAND2_365(G1273,G1102,G1198);
  nand NAND2_366(G1274,G24,G1201);
  nand NAND2_367(G1275,G1105,G1201);
  nand NAND2_368(G1276,G25,G1204);
  nand NAND2_369(G1277,G1108,G1204);
  nand NAND2_370(G1278,G26,G1207);
  nand NAND2_371(G1279,G1111,G1207);
  nand NAND2_372(G1280,G27,G1210);
  nand NAND2_373(G1281,G1114,G1210);
  nand NAND2_374(G1282,G28,G1213);
  nand NAND2_375(G1283,G1117,G1213);
  nand NAND2_376(G1284,G29,G1216);
  nand NAND2_377(G1285,G1120,G1216);
  nand NAND2_378(G1286,G30,G1219);
  nand NAND2_379(G1287,G1123,G1219);
  nand NAND2_380(G1288,G31,G1222);
  nand NAND2_381(G1289,G1126,G1222);
  nand NAND2_382(G1290,G32,G1225);
  nand NAND2_383(G1291,G1129,G1225);
  nand NAND2_384(G1292,G1228,G1229);
  nand NAND2_385(G1293,G1230,G1231);
  nand NAND2_386(G1294,G1232,G1233);
  nand NAND2_387(G1295,G1234,G1235);
  nand NAND2_388(G1296,G1236,G1237);
  nand NAND2_389(G1297,G1238,G1239);
  nand NAND2_390(G1298,G1240,G1241);
  nand NAND2_391(G1299,G1242,G1243);
  nand NAND2_392(G1300,G1244,G1245);
  nand NAND2_393(G1301,G1246,G1247);
  nand NAND2_394(G1302,G1248,G1249);
  nand NAND2_395(G1303,G1250,G1251);
  nand NAND2_396(G1304,G1252,G1253);
  nand NAND2_397(G1305,G1254,G1255);
  nand NAND2_398(G1306,G1256,G1257);
  nand NAND2_399(G1307,G1258,G1259);
  nand NAND2_400(G1308,G1260,G1261);
  nand NAND2_401(G1309,G1262,G1263);
  nand NAND2_402(G1310,G1264,G1265);
  nand NAND2_403(G1311,G1266,G1267);
  nand NAND2_404(G1312,G1268,G1269);
  nand NAND2_405(G1313,G1270,G1271);
  nand NAND2_406(G1314,G1272,G1273);
  nand NAND2_407(G1315,G1274,G1275);
  nand NAND2_408(G1316,G1276,G1277);
  nand NAND2_409(G1317,G1278,G1279);
  nand NAND2_410(G1318,G1280,G1281);
  nand NAND2_411(G1319,G1282,G1283);
  nand NAND2_412(G1320,G1284,G1285);
  nand NAND2_413(G1321,G1286,G1287);
  nand NAND2_414(G1322,G1288,G1289);
  nand NAND2_415(G1323,G1290,G1291);
  not NOT_40(G1324,G1292);
  not NOT_41(G1325,G1293);
  not NOT_42(G1326,G1294);
  not NOT_43(G1327,G1295);
  not NOT_44(G1328,G1296);
  not NOT_45(G1329,G1297);
  not NOT_46(G1330,G1298);
  not NOT_47(G1331,G1299);
  not NOT_48(G1332,G1300);
  not NOT_49(G1333,G1301);
  not NOT_50(G1334,G1302);
  not NOT_51(G1335,G1303);
  not NOT_52(G1336,G1304);
  not NOT_53(G1337,G1305);
  not NOT_54(G1338,G1306);
  not NOT_55(G1339,G1307);
  not NOT_56(G1340,G1308);
  not NOT_57(G1341,G1309);
  not NOT_58(G1342,G1310);
  not NOT_59(G1343,G1311);
  not NOT_60(G1344,G1312);
  not NOT_61(G1345,G1313);
  not NOT_62(G1346,G1314);
  not NOT_63(G1347,G1315);
  not NOT_64(G1348,G1316);
  not NOT_65(G1349,G1317);
  not NOT_66(G1350,G1318);
  not NOT_67(G1351,G1319);
  not NOT_68(G1352,G1320);
  not NOT_69(G1353,G1321);
  not NOT_70(G1354,G1322);
  not NOT_71(G1355,G1323);

endmodule

