
module c880 ( N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, 
        N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, 
        N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, 
        N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, 
        N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, 
        N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, 
        N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31 );
  input N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73,
         N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106,
         N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152,
         N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207,
         N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268,
         keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5,
         keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11,
         keyinput12, keyinput13, keyinput14, keyinput15, keyinput16,
         keyinput17, keyinput18, keyinput19, keyinput20, keyinput21,
         keyinput22, keyinput23, keyinput24, keyinput25, keyinput26,
         keyinput27, keyinput28, keyinput29, keyinput30, keyinput31;
  output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446,
         N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866,
         N874, N878, N879, N880;
  wire   n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  XNOR2X1 U227 ( .IN1(n214), .IN2(keyinput30), .Q(N880) );
  NAND3X0 U228 ( .IN1(n215), .IN2(n216), .IN3(n217), .QN(n214) );
  OA222X1 U229 ( .IN1(n218), .IN2(n219), .IN3(n220), .IN4(n221), .IN5(n222), 
        .IN6(n223), .Q(n217) );
  XOR2X1 U230 ( .IN1(keyinput26), .IN2(n224), .Q(n221) );
  OA22X1 U231 ( .IN1(n225), .IN2(n226), .IN3(n227), .IN4(n228), .Q(n224) );
  NAND2X0 U232 ( .IN1(n229), .IN2(n230), .QN(n226) );
  OA21X1 U233 ( .IN1(n231), .IN2(n232), .IN3(n227), .Q(n225) );
  INVX0 U234 ( .INP(n233), .ZN(n227) );
  NAND2X0 U235 ( .IN1(N96), .IN2(N210), .QN(n216) );
  MUX21X1 U236 ( .IN1(n234), .IN2(n235), .S(n232), .Q(n215) );
  INVX0 U237 ( .INP(n228), .ZN(n232) );
  NAND2X0 U238 ( .IN1(N228), .IN2(n236), .QN(n234) );
  NAND4X0 U239 ( .IN1(n237), .IN2(n238), .IN3(n239), .IN4(n240), .QN(N879) );
  AOI222X1 U240 ( .IN1(n241), .IN2(N165), .IN3(n242), .IN4(N237), .IN5(n243), 
        .IN6(N246), .QN(n240) );
  XOR2X1 U241 ( .IN1(n244), .IN2(keyinput29), .Q(n239) );
  NAND2X0 U242 ( .IN1(n245), .IN2(N219), .QN(n244) );
  XOR2X1 U243 ( .IN1(n246), .IN2(n247), .Q(n245) );
  NAND3X0 U244 ( .IN1(n229), .IN2(n230), .IN3(n228), .QN(n246) );
  NAND2X0 U245 ( .IN1(N91), .IN2(N210), .QN(n238) );
  XOR2X1 U246 ( .IN1(keyinput21), .IN2(n248), .Q(n237) );
  AND2X1 U247 ( .IN1(N228), .IN2(n247), .Q(n248) );
  NOR2X0 U248 ( .IN1(n242), .IN2(n249), .QN(n247) );
  XOR2X1 U249 ( .IN1(keyinput31), .IN2(n250), .Q(N878) );
  NOR2X0 U250 ( .IN1(n251), .IN2(n252), .QN(n250) );
  AO221X1 U251 ( .IN1(N159), .IN2(n241), .IN3(N268), .IN4(N210), .IN5(n253), 
        .Q(n252) );
  XOR2X1 U252 ( .IN1(keyinput20), .IN2(n254), .Q(n253) );
  NOR2X0 U253 ( .IN1(n255), .IN2(n256), .QN(n254) );
  AO222X1 U254 ( .IN1(n257), .IN2(N237), .IN3(n258), .IN4(N219), .IN5(N246), 
        .IN6(n259), .Q(n251) );
  XNOR2X1 U255 ( .IN1(n256), .IN2(n260), .Q(n258) );
  AO21X1 U256 ( .IN1(n261), .IN2(n262), .IN3(n257), .Q(n256) );
  NAND3X0 U257 ( .IN1(n263), .IN2(n264), .IN3(n265), .QN(N874) );
  AOI222X1 U258 ( .IN1(N177), .IN2(n241), .IN3(n266), .IN4(N219), .IN5(n267), 
        .IN6(N246), .QN(n265) );
  OAI22X1 U259 ( .IN1(n268), .IN2(n269), .IN3(n270), .IN4(n233), .QN(n266) );
  NAND2X0 U260 ( .IN1(n271), .IN2(n272), .QN(n233) );
  OA21X1 U261 ( .IN1(n273), .IN2(n274), .IN3(n275), .Q(n269) );
  NOR2X0 U262 ( .IN1(n276), .IN2(n272), .QN(n268) );
  NAND2X0 U263 ( .IN1(N210), .IN2(N101), .QN(n264) );
  XOR2X1 U264 ( .IN1(keyinput23), .IN2(n277), .Q(n263) );
  MUX21X1 U265 ( .IN1(N237), .IN2(n278), .S(n271), .Q(n277) );
  NOR2X0 U266 ( .IN1(n270), .IN2(n255), .QN(n278) );
  AO21X1 U267 ( .IN1(n279), .IN2(n260), .IN3(n257), .Q(N866) );
  NOR2X0 U268 ( .IN1(n262), .IN2(n261), .QN(n257) );
  OAI221X1 U269 ( .IN1(n249), .IN2(n228), .IN3(n280), .IN4(n249), .IN5(n281), 
        .QN(n260) );
  INVX0 U270 ( .INP(n242), .ZN(n281) );
  XNOR2X1 U271 ( .IN1(n282), .IN2(keyinput16), .Q(n242) );
  NAND2X0 U272 ( .IN1(N165), .IN2(n243), .QN(n282) );
  AND2X1 U273 ( .IN1(n230), .IN2(n229), .Q(n280) );
  OR2X1 U274 ( .IN1(n272), .IN2(n231), .Q(n229) );
  INVX0 U275 ( .INP(n236), .ZN(n231) );
  AO21X1 U276 ( .IN1(n275), .IN2(n283), .IN3(n270), .Q(n272) );
  NOR2X0 U277 ( .IN1(n267), .IN2(N177), .QN(n270) );
  OR2X1 U278 ( .IN1(n274), .IN2(n273), .Q(n283) );
  NAND2X0 U279 ( .IN1(n276), .IN2(n236), .QN(n230) );
  NAND2X0 U280 ( .IN1(n222), .IN2(n218), .QN(n236) );
  INVX0 U281 ( .INP(n284), .ZN(n222) );
  INVX0 U282 ( .INP(n271), .ZN(n276) );
  NAND2X0 U283 ( .IN1(N177), .IN2(n267), .QN(n271) );
  AO222X1 U284 ( .IN1(N152), .IN2(N138), .IN3(n285), .IN4(n286), .IN5(N106), 
        .IN6(n287), .Q(n267) );
  NAND2X0 U285 ( .IN1(n288), .IN2(n289), .QN(n286) );
  INVX0 U286 ( .INP(N153), .ZN(n289) );
  NAND2X0 U287 ( .IN1(N171), .IN2(n284), .QN(n228) );
  AO222X1 U288 ( .IN1(N101), .IN2(n287), .IN3(n290), .IN4(n285), .IN5(N138), 
        .IN6(N17), .Q(n284) );
  NAND2X0 U289 ( .IN1(n291), .IN2(n288), .QN(n290) );
  INVX0 U290 ( .INP(N149), .ZN(n291) );
  NOR2X0 U291 ( .IN1(n243), .IN2(N165), .QN(n249) );
  AO222X1 U292 ( .IN1(N96), .IN2(n287), .IN3(n292), .IN4(n285), .IN5(N138), 
        .IN6(N51), .Q(n243) );
  NAND2X0 U293 ( .IN1(n293), .IN2(n288), .QN(n285) );
  NAND2X0 U294 ( .IN1(n294), .IN2(n288), .QN(n292) );
  INVX0 U295 ( .INP(N146), .ZN(n294) );
  NAND2X0 U296 ( .IN1(n261), .IN2(n262), .QN(n279) );
  INVX0 U297 ( .INP(N159), .ZN(n262) );
  INVX0 U298 ( .INP(n259), .ZN(n261) );
  AO221X1 U299 ( .IN1(n295), .IN2(N143), .IN3(N91), .IN4(n287), .IN5(n296), 
        .Q(n259) );
  AO21X1 U300 ( .IN1(N8), .IN2(N138), .IN3(n297), .Q(n296) );
  XOR2X1 U301 ( .IN1(n288), .IN2(keyinput8), .Q(n297) );
  NAND2X0 U302 ( .IN1(N17), .IN2(n298), .QN(n288) );
  INVX0 U303 ( .INP(n293), .ZN(n295) );
  NAND3X0 U304 ( .IN1(N447), .IN2(n299), .IN3(N55), .QN(n293) );
  NAND3X0 U305 ( .IN1(n300), .IN2(n301), .IN3(n302), .QN(N863) );
  OA222X1 U306 ( .IN1(n255), .IN2(n303), .IN3(n304), .IN4(n220), .IN5(n275), 
        .IN6(n235), .Q(n302) );
  XOR2X1 U307 ( .IN1(n305), .IN2(keyinput18), .Q(n275) );
  NAND2X0 U308 ( .IN1(N183), .IN2(n306), .QN(n305) );
  XNOR2X1 U309 ( .IN1(n303), .IN2(n273), .Q(n304) );
  XNOR2X1 U310 ( .IN1(keyinput24), .IN2(n307), .Q(n273) );
  OA221X1 U311 ( .IN1(n308), .IN2(n309), .IN3(n309), .IN4(n310), .IN5(n311), 
        .Q(n307) );
  XNOR2X1 U312 ( .IN1(n312), .IN2(keyinput22), .Q(n311) );
  AND2X1 U313 ( .IN1(n313), .IN2(n314), .Q(n308) );
  AO21X1 U314 ( .IN1(N183), .IN2(n306), .IN3(n274), .Q(n303) );
  XOR2X1 U315 ( .IN1(n315), .IN2(keyinput17), .Q(n274) );
  NAND2X0 U316 ( .IN1(n316), .IN2(n317), .QN(n315) );
  XOR2X1 U317 ( .IN1(n318), .IN2(keyinput3), .Q(n301) );
  NAND2X0 U318 ( .IN1(N210), .IN2(N106), .QN(n318) );
  OA22X1 U319 ( .IN1(n316), .IN2(n223), .IN3(n317), .IN4(n219), .Q(n300) );
  INVX0 U320 ( .INP(N246), .ZN(n223) );
  INVX0 U321 ( .INP(n306), .ZN(n316) );
  AO221X1 U322 ( .IN1(N111), .IN2(n287), .IN3(N143), .IN4(n319), .IN5(n320), 
        .Q(n306) );
  NAND3X0 U323 ( .IN1(n321), .IN2(n322), .IN3(n323), .QN(N850) );
  OA222X1 U324 ( .IN1(n324), .IN2(n235), .IN3(n325), .IN4(n220), .IN5(n255), 
        .IN6(n326), .Q(n323) );
  INVX0 U325 ( .INP(N228), .ZN(n255) );
  INVX0 U326 ( .INP(N219), .ZN(n220) );
  XOR2X1 U327 ( .IN1(n326), .IN2(N261), .Q(n325) );
  OAI21X1 U328 ( .IN1(n327), .IN2(N201), .IN3(n324), .QN(n326) );
  INVX0 U329 ( .INP(N237), .ZN(n235) );
  XOR2X1 U330 ( .IN1(n328), .IN2(keyinput19), .Q(n322) );
  AO22X1 U331 ( .IN1(N267), .IN2(N255), .IN3(N246), .IN4(n327), .Q(n328) );
  AOI22X1 U332 ( .IN1(N201), .IN2(n241), .IN3(N121), .IN4(N210), .QN(n321) );
  XOR3X1 U333 ( .IN1(N207), .IN2(n329), .IN3(n330), .Q(N768) );
  NOR3X0 U334 ( .IN1(n331), .IN2(keyinput15), .IN3(n332), .QN(n330) );
  NOR2X0 U335 ( .IN1(n333), .IN2(n334), .QN(n332) );
  XOR2X1 U336 ( .IN1(n335), .IN2(keyinput12), .Q(n331) );
  NAND2X0 U337 ( .IN1(n333), .IN2(n334), .QN(n335) );
  XOR3X1 U338 ( .IN1(N165), .IN2(N159), .IN3(n336), .Q(n333) );
  XOR2X1 U339 ( .IN1(n218), .IN2(N177), .Q(n336) );
  INVX0 U340 ( .INP(N171), .ZN(n218) );
  OA22X1 U341 ( .IN1(n337), .IN2(n338), .IN3(n339), .IN4(n340), .Q(n329) );
  MUX21X1 U342 ( .IN1(n341), .IN2(n342), .S(n343), .Q(n340) );
  AND2X1 U343 ( .IN1(n342), .IN2(n343), .Q(n337) );
  XNOR2X1 U344 ( .IN1(n317), .IN2(N189), .Q(n343) );
  INVX0 U345 ( .INP(N183), .ZN(n317) );
  OAI21X1 U346 ( .IN1(n339), .IN2(n338), .IN3(n341), .QN(n342) );
  INVX0 U347 ( .INP(keyinput5), .ZN(n341) );
  XOR2X1 U348 ( .IN1(N195), .IN2(N201), .Q(n338) );
  INVX0 U349 ( .INP(keyinput6), .ZN(n339) );
  XOR3X1 U350 ( .IN1(N121), .IN2(n344), .IN3(n345), .Q(N767) );
  XOR3X1 U351 ( .IN1(N116), .IN2(N111), .IN3(n346), .Q(n345) );
  NOR2X0 U352 ( .IN1(n347), .IN2(n348), .QN(n346) );
  XOR2X1 U353 ( .IN1(n349), .IN2(keyinput10), .Q(n348) );
  NAND2X0 U354 ( .IN1(n350), .IN2(n334), .QN(n349) );
  XOR2X1 U355 ( .IN1(n351), .IN2(keyinput9), .Q(n347) );
  OR2X1 U356 ( .IN1(n350), .IN2(n334), .Q(n351) );
  INVX0 U357 ( .INP(N130), .ZN(n334) );
  AO21X1 U358 ( .IN1(n352), .IN2(n353), .IN3(n354), .Q(n350) );
  XOR2X1 U359 ( .IN1(n355), .IN2(keyinput7), .Q(n354) );
  NAND2X0 U360 ( .IN1(n356), .IN2(n357), .QN(n355) );
  XOR2X1 U361 ( .IN1(N96), .IN2(N91), .Q(n357) );
  INVX0 U362 ( .INP(n353), .ZN(n356) );
  AO21X1 U363 ( .IN1(n358), .IN2(n359), .IN3(n360), .Q(n353) );
  XOR2X1 U364 ( .IN1(keyinput2), .IN2(n361), .Q(n360) );
  NOR2X0 U365 ( .IN1(n359), .IN2(n358), .QN(n361) );
  INVX0 U366 ( .INP(N106), .ZN(n359) );
  INVX0 U367 ( .INP(N101), .ZN(n358) );
  XNOR2X1 U368 ( .IN1(N91), .IN2(N96), .Q(n352) );
  XOR2X1 U369 ( .IN1(N135), .IN2(N126), .Q(n344) );
  AND4X1 U370 ( .IN1(n362), .IN2(n363), .IN3(N59), .IN4(N55), .Q(N449) );
  AND2X1 U371 ( .IN1(N74), .IN2(N68), .Q(n362) );
  AND3X1 U372 ( .IN1(n363), .IN2(N55), .IN3(n364), .Q(N448) );
  XOR2X1 U373 ( .IN1(n365), .IN2(keyinput1), .Q(n364) );
  NAND2X0 U374 ( .IN1(N68), .IN2(N29), .QN(n365) );
  NAND2X0 U375 ( .IN1(N36), .IN2(n366), .QN(N422) );
  NAND3X0 U376 ( .IN1(N59), .IN2(N80), .IN3(N36), .QN(N421) );
  NAND3X0 U377 ( .IN1(N80), .IN2(N75), .IN3(N59), .QN(N420) );
  NAND2X0 U378 ( .IN1(n367), .IN2(n368), .QN(N446) );
  XOR2X1 U379 ( .IN1(n369), .IN2(keyinput0), .Q(n367) );
  AND2X1 U380 ( .IN1(N90), .IN2(n370), .Q(N423) );
  NAND2X0 U381 ( .IN1(n368), .IN2(n371), .QN(N419) );
  XOR2X1 U382 ( .IN1(keyinput0), .IN2(N390), .Q(n371) );
  AND4X1 U383 ( .IN1(N13), .IN2(N17), .IN3(N26), .IN4(N1), .Q(n368) );
  AND2X1 U384 ( .IN1(N86), .IN2(N85), .Q(N391) );
  INVX0 U385 ( .INP(n369), .ZN(N390) );
  NAND3X0 U386 ( .IN1(N42), .IN2(N29), .IN3(N36), .QN(n369) );
  AND3X1 U387 ( .IN1(N80), .IN2(N29), .IN3(N36), .Q(N389) );
  AND3X1 U388 ( .IN1(N75), .IN2(N29), .IN3(N42), .Q(N388) );
  AND2X1 U389 ( .IN1(N89), .IN2(n370), .Q(N450) );
  OR2X1 U390 ( .IN1(N87), .IN2(N88), .Q(n370) );
  XOR2X1 U391 ( .IN1(keyinput28), .IN2(n372), .Q(N865) );
  NOR2X0 U392 ( .IN1(n373), .IN2(n374), .QN(n372) );
  AO222X1 U393 ( .IN1(N210), .IN2(N116), .IN3(n241), .IN4(N195), .IN5(N260), 
        .IN6(N255), .Q(n374) );
  AO221X1 U394 ( .IN1(n375), .IN2(N219), .IN3(n376), .IN4(N228), .IN5(n377), 
        .Q(n373) );
  AO22X1 U395 ( .IN1(N246), .IN2(n378), .IN3(N237), .IN4(n379), .Q(n377) );
  INVX0 U396 ( .INP(n310), .ZN(n379) );
  INVX0 U397 ( .INP(n380), .ZN(n376) );
  MUX21X1 U398 ( .IN1(n381), .IN2(n382), .S(keyinput25), .Q(n375) );
  XOR2X1 U399 ( .IN1(n383), .IN2(n380), .Q(n382) );
  NOR2X0 U400 ( .IN1(n383), .IN2(n380), .QN(n381) );
  NAND2X0 U401 ( .IN1(n310), .IN2(n384), .QN(n380) );
  NOR2X0 U402 ( .IN1(n385), .IN2(n386), .QN(n383) );
  XOR2X1 U403 ( .IN1(keyinput27), .IN2(n387), .Q(N864) );
  NOR2X0 U404 ( .IN1(n388), .IN2(n389), .QN(n387) );
  AO222X1 U405 ( .IN1(N210), .IN2(N111), .IN3(n241), .IN4(N189), .IN5(N259), 
        .IN6(N255), .Q(n389) );
  INVX0 U406 ( .INP(n219), .ZN(n241) );
  NAND4X0 U407 ( .IN1(n366), .IN2(N55), .IN3(n363), .IN4(n390), .QN(n219) );
  AND3X1 U408 ( .IN1(N72), .IN2(N68), .IN3(N73), .Q(n390) );
  AO221X1 U409 ( .IN1(n391), .IN2(N219), .IN3(n392), .IN4(N228), .IN5(n393), 
        .Q(n388) );
  AO22X1 U410 ( .IN1(N246), .IN2(n394), .IN3(N237), .IN4(n312), .Q(n393) );
  XOR2X1 U411 ( .IN1(n395), .IN2(n392), .Q(n391) );
  NOR2X0 U412 ( .IN1(n312), .IN2(n309), .QN(n392) );
  NOR2X0 U413 ( .IN1(n394), .IN2(N189), .QN(n309) );
  AND2X1 U414 ( .IN1(N189), .IN2(n394), .Q(n312) );
  XOR2X1 U415 ( .IN1(n396), .IN2(keyinput13), .Q(n394) );
  AO221X1 U416 ( .IN1(N116), .IN2(n287), .IN3(N146), .IN4(n319), .IN5(n320), 
        .Q(n396) );
  NAND3X0 U417 ( .IN1(n313), .IN2(n310), .IN3(n314), .QN(n395) );
  NAND2X0 U418 ( .IN1(n386), .IN2(n384), .QN(n314) );
  INVX0 U419 ( .INP(n324), .ZN(n386) );
  NAND2X0 U420 ( .IN1(N201), .IN2(n327), .QN(n324) );
  NAND2X0 U421 ( .IN1(N195), .IN2(n378), .QN(n310) );
  NAND2X0 U422 ( .IN1(n385), .IN2(n384), .QN(n313) );
  OR2X1 U423 ( .IN1(n378), .IN2(N195), .Q(n384) );
  XNOR2X1 U424 ( .IN1(n397), .IN2(keyinput14), .Q(n378) );
  AO221X1 U425 ( .IN1(N121), .IN2(n287), .IN3(N149), .IN4(n319), .IN5(n320), 
        .Q(n397) );
  INVX0 U426 ( .INP(n398), .ZN(n320) );
  OA21X1 U427 ( .IN1(n327), .IN2(N201), .IN3(N261), .Q(n385) );
  NAND3X0 U428 ( .IN1(n399), .IN2(n398), .IN3(n400), .QN(n327) );
  XOR2X1 U429 ( .IN1(n401), .IN2(keyinput11), .Q(n400) );
  NAND2X0 U430 ( .IN1(N126), .IN2(n287), .QN(n401) );
  AO22X1 U431 ( .IN1(n402), .IN2(n403), .IN3(n404), .IN4(n405), .Q(n287) );
  INVX0 U432 ( .INP(n299), .ZN(n405) );
  NOR2X0 U433 ( .IN1(n406), .IN2(n407), .QN(n404) );
  XNOR2X1 U434 ( .IN1(N42), .IN2(N17), .Q(n406) );
  NAND2X0 U435 ( .IN1(n366), .IN2(N75), .QN(n403) );
  AND2X1 U436 ( .IN1(N42), .IN2(N59), .Q(n366) );
  XNOR2X1 U437 ( .IN1(n408), .IN2(keyinput4), .Q(n402) );
  NAND4X0 U438 ( .IN1(N8), .IN2(N17), .IN3(N51), .IN4(N1), .QN(n408) );
  NAND2X0 U439 ( .IN1(N55), .IN2(n298), .QN(n398) );
  AND4X1 U440 ( .IN1(N447), .IN2(n409), .IN3(N29), .IN4(n410), .Q(n298) );
  AND2X1 U441 ( .IN1(N75), .IN2(N80), .Q(n410) );
  INVX0 U442 ( .INP(N268), .ZN(n409) );
  NAND2X0 U443 ( .IN1(N153), .IN2(n319), .QN(n399) );
  NAND2X0 U444 ( .IN1(N1), .IN2(n411), .QN(n319) );
  NAND3X0 U445 ( .IN1(N447), .IN2(n299), .IN3(N17), .QN(n411) );
  NAND2X0 U446 ( .IN1(N59), .IN2(N156), .QN(n299) );
  INVX0 U447 ( .INP(n407), .ZN(N447) );
  NAND3X0 U448 ( .IN1(N26), .IN2(N1), .IN3(N51), .QN(n407) );
  AND2X1 U449 ( .IN1(N17), .IN2(n363), .Q(N418) );
  AND3X1 U450 ( .IN1(N8), .IN2(N1), .IN3(N13), .Q(n363) );
endmodule

