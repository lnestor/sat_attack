
module c6288 ( N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, 
        N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, 
        N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, N1901, 
        N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, 
        N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, 
        N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31 );
  input N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205,
         N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392,
         N409, N426, N443, N460, N477, N494, N511, N528, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31;
  output N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241,
         N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180,
         N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280,
         N6287, N6288;
  wire   n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927;

  NAND2X0 U1526 ( .IN1(n1495), .IN2(n1496), .QN(N6288) );
  NAND3X0 U1527 ( .IN1(n1497), .IN2(n1498), .IN3(n1499), .QN(n1496) );
  NOR2X0 U1528 ( .IN1(n1500), .IN2(n1501), .QN(N6287) );
  OA21X1 U1529 ( .IN1(n1502), .IN2(n1503), .IN3(n1504), .Q(n1501) );
  INVX0 U1530 ( .INP(N528), .ZN(n1503) );
  INVX0 U1531 ( .INP(n1495), .ZN(n1500) );
  AO21X1 U1532 ( .IN1(n1497), .IN2(n1498), .IN3(n1499), .Q(n1495) );
  XNOR2X1 U1533 ( .IN1(n1505), .IN2(n1504), .Q(n1499) );
  NAND2X0 U1534 ( .IN1(n1506), .IN2(n1507), .QN(n1504) );
  AO21X1 U1535 ( .IN1(N256), .IN2(N511), .IN3(n1508), .Q(n1506) );
  NAND2X0 U1536 ( .IN1(N528), .IN2(N256), .QN(n1505) );
  NAND2X0 U1537 ( .IN1(n1497), .IN2(n1509), .QN(N6280) );
  NAND3X0 U1538 ( .IN1(n1510), .IN2(n1511), .IN3(n1512), .QN(n1509) );
  AO21X1 U1539 ( .IN1(n1510), .IN2(n1511), .IN3(n1512), .Q(n1497) );
  NAND2X0 U1540 ( .IN1(n1498), .IN2(n1513), .QN(n1512) );
  NAND3X0 U1541 ( .IN1(n1514), .IN2(n1515), .IN3(n1516), .QN(n1513) );
  AO21X1 U1542 ( .IN1(n1514), .IN2(n1515), .IN3(n1516), .Q(n1498) );
  NAND2X0 U1543 ( .IN1(n1507), .IN2(n1517), .QN(n1516) );
  NAND3X0 U1544 ( .IN1(n1518), .IN2(N239), .IN3(N528), .QN(n1517) );
  AO21X1 U1545 ( .IN1(N528), .IN2(N239), .IN3(n1518), .Q(n1507) );
  XNOR2X1 U1546 ( .IN1(n1508), .IN2(n1519), .Q(n1518) );
  AND2X1 U1547 ( .IN1(N511), .IN2(N256), .Q(n1519) );
  AND2X1 U1548 ( .IN1(n1520), .IN2(n1521), .Q(n1508) );
  AO21X1 U1549 ( .IN1(N256), .IN2(N494), .IN3(n1522), .Q(n1520) );
  INVX0 U1550 ( .INP(n1523), .ZN(n1511) );
  NAND2X0 U1551 ( .IN1(n1510), .IN2(n1524), .QN(N6270) );
  NAND3X0 U1552 ( .IN1(n1525), .IN2(n1526), .IN3(n1527), .QN(n1524) );
  AO21X1 U1553 ( .IN1(n1525), .IN2(n1526), .IN3(n1527), .Q(n1510) );
  AO21X1 U1554 ( .IN1(n1528), .IN2(n1529), .IN3(n1523), .Q(n1527) );
  NOR2X0 U1555 ( .IN1(n1529), .IN2(n1528), .QN(n1523) );
  NAND2X0 U1556 ( .IN1(n1514), .IN2(n1530), .QN(n1529) );
  NAND3X0 U1557 ( .IN1(N528), .IN2(n1531), .IN3(N222), .QN(n1530) );
  AO21X1 U1558 ( .IN1(N222), .IN2(N528), .IN3(n1531), .Q(n1514) );
  NAND2X0 U1559 ( .IN1(n1515), .IN2(n1532), .QN(n1531) );
  NAND3X0 U1560 ( .IN1(n1533), .IN2(n1534), .IN3(n1535), .QN(n1532) );
  AO21X1 U1561 ( .IN1(n1533), .IN2(n1534), .IN3(n1535), .Q(n1515) );
  NAND2X0 U1562 ( .IN1(n1521), .IN2(n1536), .QN(n1535) );
  NAND3X0 U1563 ( .IN1(N511), .IN2(N239), .IN3(n1537), .QN(n1536) );
  AO21X1 U1564 ( .IN1(N511), .IN2(N239), .IN3(n1537), .Q(n1521) );
  XNOR2X1 U1565 ( .IN1(n1522), .IN2(n1538), .Q(n1537) );
  AND2X1 U1566 ( .IN1(N494), .IN2(N256), .Q(n1538) );
  AND2X1 U1567 ( .IN1(n1539), .IN2(n1540), .Q(n1522) );
  AO21X1 U1568 ( .IN1(N256), .IN2(N477), .IN3(n1541), .Q(n1539) );
  XNOR2X1 U1569 ( .IN1(keyinput26), .IN2(n1542), .Q(n1528) );
  OA21X1 U1570 ( .IN1(n1543), .IN2(n1544), .IN3(n1545), .Q(n1542) );
  NAND2X0 U1571 ( .IN1(n1525), .IN2(n1546), .QN(N6260) );
  NAND3X0 U1572 ( .IN1(n1547), .IN2(n1548), .IN3(n1549), .QN(n1546) );
  AO21X1 U1573 ( .IN1(n1547), .IN2(n1548), .IN3(n1549), .Q(n1525) );
  NAND2X0 U1574 ( .IN1(n1526), .IN2(n1550), .QN(n1549) );
  NAND3X0 U1575 ( .IN1(n1551), .IN2(n1552), .IN3(n1553), .QN(n1550) );
  AO21X1 U1576 ( .IN1(n1551), .IN2(n1552), .IN3(n1553), .Q(n1526) );
  NAND2X0 U1577 ( .IN1(n1545), .IN2(n1554), .QN(n1553) );
  NAND3X0 U1578 ( .IN1(N528), .IN2(n1555), .IN3(N205), .QN(n1554) );
  AO21X1 U1579 ( .IN1(N205), .IN2(N528), .IN3(n1555), .Q(n1545) );
  XNOR2X1 U1580 ( .IN1(n1543), .IN2(n1544), .Q(n1555) );
  AND2X1 U1581 ( .IN1(n1556), .IN2(n1557), .Q(n1544) );
  NAND2X0 U1582 ( .IN1(n1533), .IN2(n1558), .QN(n1543) );
  NAND3X0 U1583 ( .IN1(N511), .IN2(n1559), .IN3(N222), .QN(n1558) );
  AO21X1 U1584 ( .IN1(N222), .IN2(N511), .IN3(n1559), .Q(n1533) );
  NAND2X0 U1585 ( .IN1(n1534), .IN2(n1560), .QN(n1559) );
  NAND3X0 U1586 ( .IN1(n1561), .IN2(n1562), .IN3(n1563), .QN(n1560) );
  AO21X1 U1587 ( .IN1(n1561), .IN2(n1562), .IN3(n1563), .Q(n1534) );
  NAND2X0 U1588 ( .IN1(n1540), .IN2(n1564), .QN(n1563) );
  NAND3X0 U1589 ( .IN1(N494), .IN2(N239), .IN3(n1565), .QN(n1564) );
  AO21X1 U1590 ( .IN1(N494), .IN2(N239), .IN3(n1565), .Q(n1540) );
  XNOR2X1 U1591 ( .IN1(n1541), .IN2(n1566), .Q(n1565) );
  AND2X1 U1592 ( .IN1(N477), .IN2(N256), .Q(n1566) );
  AND2X1 U1593 ( .IN1(n1567), .IN2(n1568), .Q(n1541) );
  AO21X1 U1594 ( .IN1(N256), .IN2(N460), .IN3(n1569), .Q(n1567) );
  NAND2X0 U1595 ( .IN1(n1547), .IN2(n1570), .QN(N6250) );
  NAND3X0 U1596 ( .IN1(n1571), .IN2(n1572), .IN3(n1573), .QN(n1570) );
  AO21X1 U1597 ( .IN1(n1571), .IN2(n1572), .IN3(n1573), .Q(n1547) );
  NAND2X0 U1598 ( .IN1(n1548), .IN2(n1574), .QN(n1573) );
  NAND3X0 U1599 ( .IN1(n1575), .IN2(n1576), .IN3(n1577), .QN(n1574) );
  AO21X1 U1600 ( .IN1(n1575), .IN2(n1576), .IN3(n1577), .Q(n1548) );
  NAND2X0 U1601 ( .IN1(n1551), .IN2(n1578), .QN(n1577) );
  NAND3X0 U1602 ( .IN1(N528), .IN2(n1579), .IN3(N188), .QN(n1578) );
  AO21X1 U1603 ( .IN1(N188), .IN2(N528), .IN3(n1579), .Q(n1551) );
  NAND2X0 U1604 ( .IN1(n1552), .IN2(n1580), .QN(n1579) );
  NAND3X0 U1605 ( .IN1(n1581), .IN2(n1582), .IN3(n1583), .QN(n1580) );
  AO21X1 U1606 ( .IN1(n1581), .IN2(n1582), .IN3(n1583), .Q(n1552) );
  NAND2X0 U1607 ( .IN1(n1557), .IN2(n1584), .QN(n1583) );
  NAND3X0 U1608 ( .IN1(N511), .IN2(n1585), .IN3(N205), .QN(n1584) );
  AO21X1 U1609 ( .IN1(N205), .IN2(N511), .IN3(n1585), .Q(n1557) );
  NAND2X0 U1610 ( .IN1(n1556), .IN2(n1586), .QN(n1585) );
  NAND4X0 U1611 ( .IN1(n1587), .IN2(n1588), .IN3(n1589), .IN4(n1590), .QN(
        n1586) );
  AO22X1 U1612 ( .IN1(n1587), .IN2(n1588), .IN3(n1589), .IN4(n1590), .Q(n1556)
         );
  NAND2X0 U1613 ( .IN1(n1591), .IN2(n1561), .QN(n1588) );
  XNOR2X1 U1614 ( .IN1(n1592), .IN2(keyinput20), .Q(n1587) );
  NAND2X0 U1615 ( .IN1(n1561), .IN2(n1593), .QN(n1592) );
  NAND2X0 U1616 ( .IN1(n1591), .IN2(n1593), .QN(n1561) );
  NAND2X0 U1617 ( .IN1(N222), .IN2(N494), .QN(n1593) );
  AND2X1 U1618 ( .IN1(n1562), .IN2(n1594), .Q(n1591) );
  NAND3X0 U1619 ( .IN1(n1595), .IN2(n1596), .IN3(n1597), .QN(n1594) );
  AO21X1 U1620 ( .IN1(n1597), .IN2(n1596), .IN3(n1595), .Q(n1562) );
  NAND2X0 U1621 ( .IN1(n1568), .IN2(n1598), .QN(n1595) );
  NAND3X0 U1622 ( .IN1(N477), .IN2(N239), .IN3(n1599), .QN(n1598) );
  AO21X1 U1623 ( .IN1(N477), .IN2(N239), .IN3(n1599), .Q(n1568) );
  XNOR2X1 U1624 ( .IN1(n1569), .IN2(n1600), .Q(n1599) );
  AND2X1 U1625 ( .IN1(N460), .IN2(N256), .Q(n1600) );
  AND2X1 U1626 ( .IN1(n1601), .IN2(n1602), .Q(n1569) );
  AO21X1 U1627 ( .IN1(n1603), .IN2(n1604), .IN3(n1605), .Q(n1601) );
  NAND2X0 U1628 ( .IN1(n1571), .IN2(n1606), .QN(N6240) );
  NAND3X0 U1629 ( .IN1(n1607), .IN2(n1608), .IN3(n1609), .QN(n1606) );
  AO21X1 U1630 ( .IN1(n1607), .IN2(n1608), .IN3(n1609), .Q(n1571) );
  NAND2X0 U1631 ( .IN1(n1572), .IN2(n1610), .QN(n1609) );
  NAND3X0 U1632 ( .IN1(n1611), .IN2(n1612), .IN3(n1613), .QN(n1610) );
  AO21X1 U1633 ( .IN1(n1611), .IN2(n1612), .IN3(n1613), .Q(n1572) );
  NAND2X0 U1634 ( .IN1(n1575), .IN2(n1614), .QN(n1613) );
  NAND3X0 U1635 ( .IN1(N528), .IN2(n1615), .IN3(N171), .QN(n1614) );
  AO21X1 U1636 ( .IN1(N171), .IN2(N528), .IN3(n1615), .Q(n1575) );
  NAND2X0 U1637 ( .IN1(n1576), .IN2(n1616), .QN(n1615) );
  NAND3X0 U1638 ( .IN1(n1617), .IN2(n1618), .IN3(n1619), .QN(n1616) );
  AO21X1 U1639 ( .IN1(n1617), .IN2(n1618), .IN3(n1619), .Q(n1576) );
  XNOR2X1 U1640 ( .IN1(n1620), .IN2(keyinput25), .Q(n1619) );
  NAND2X0 U1641 ( .IN1(n1581), .IN2(n1621), .QN(n1620) );
  NAND3X0 U1642 ( .IN1(N511), .IN2(n1622), .IN3(N188), .QN(n1621) );
  AO21X1 U1643 ( .IN1(N188), .IN2(N511), .IN3(n1622), .Q(n1581) );
  NAND2X0 U1644 ( .IN1(n1582), .IN2(n1623), .QN(n1622) );
  NAND3X0 U1645 ( .IN1(n1624), .IN2(n1625), .IN3(n1626), .QN(n1623) );
  AO21X1 U1646 ( .IN1(n1624), .IN2(n1625), .IN3(n1626), .Q(n1582) );
  NAND2X0 U1647 ( .IN1(n1589), .IN2(n1627), .QN(n1626) );
  NAND3X0 U1648 ( .IN1(N494), .IN2(n1628), .IN3(N205), .QN(n1627) );
  AO21X1 U1649 ( .IN1(N205), .IN2(N494), .IN3(n1628), .Q(n1589) );
  NAND2X0 U1650 ( .IN1(n1590), .IN2(n1629), .QN(n1628) );
  NAND3X0 U1651 ( .IN1(n1630), .IN2(n1631), .IN3(n1632), .QN(n1629) );
  AO21X1 U1652 ( .IN1(n1630), .IN2(n1631), .IN3(n1632), .Q(n1590) );
  NAND2X0 U1653 ( .IN1(n1597), .IN2(n1633), .QN(n1632) );
  NAND3X0 U1654 ( .IN1(N477), .IN2(n1634), .IN3(N222), .QN(n1633) );
  XNOR2X1 U1655 ( .IN1(keyinput18), .IN2(n1635), .Q(n1597) );
  AOI21X1 U1656 ( .IN1(N477), .IN2(N222), .IN3(n1634), .QN(n1635) );
  NAND2X0 U1657 ( .IN1(n1596), .IN2(n1636), .QN(n1634) );
  NAND3X0 U1658 ( .IN1(n1637), .IN2(n1638), .IN3(n1639), .QN(n1636) );
  AO21X1 U1659 ( .IN1(n1637), .IN2(n1638), .IN3(n1639), .Q(n1596) );
  NAND2X0 U1660 ( .IN1(n1602), .IN2(n1640), .QN(n1639) );
  NAND3X0 U1661 ( .IN1(N239), .IN2(n1641), .IN3(N460), .QN(n1640) );
  AO21X1 U1662 ( .IN1(N460), .IN2(N239), .IN3(n1641), .Q(n1602) );
  XOR2X1 U1663 ( .IN1(n1642), .IN2(n1605), .Q(n1641) );
  XOR2X1 U1664 ( .IN1(n1643), .IN2(keyinput2), .Q(n1605) );
  NAND2X0 U1665 ( .IN1(N443), .IN2(N256), .QN(n1643) );
  NAND2X0 U1666 ( .IN1(n1604), .IN2(n1603), .QN(n1642) );
  NAND2X0 U1667 ( .IN1(n1607), .IN2(n1644), .QN(N6230) );
  NAND3X0 U1668 ( .IN1(n1645), .IN2(n1646), .IN3(n1647), .QN(n1644) );
  AO21X1 U1669 ( .IN1(n1645), .IN2(n1646), .IN3(n1647), .Q(n1607) );
  NAND2X0 U1670 ( .IN1(n1608), .IN2(n1648), .QN(n1647) );
  NAND3X0 U1671 ( .IN1(n1649), .IN2(n1650), .IN3(n1651), .QN(n1648) );
  AO21X1 U1672 ( .IN1(n1649), .IN2(n1650), .IN3(n1651), .Q(n1608) );
  NAND2X0 U1673 ( .IN1(n1611), .IN2(n1652), .QN(n1651) );
  NAND3X0 U1674 ( .IN1(N528), .IN2(n1653), .IN3(N154), .QN(n1652) );
  AO21X1 U1675 ( .IN1(N154), .IN2(N528), .IN3(n1653), .Q(n1611) );
  NAND2X0 U1676 ( .IN1(n1612), .IN2(n1654), .QN(n1653) );
  NAND3X0 U1677 ( .IN1(n1655), .IN2(n1656), .IN3(n1657), .QN(n1654) );
  AO21X1 U1678 ( .IN1(n1655), .IN2(n1656), .IN3(n1657), .Q(n1612) );
  OA21X1 U1679 ( .IN1(n1658), .IN2(n1659), .IN3(n1660), .Q(n1657) );
  NAND2X0 U1680 ( .IN1(n1661), .IN2(n1617), .QN(n1656) );
  XOR2X1 U1681 ( .IN1(n1662), .IN2(keyinput24), .Q(n1655) );
  NAND2X0 U1682 ( .IN1(n1617), .IN2(n1663), .QN(n1662) );
  NAND2X0 U1683 ( .IN1(n1661), .IN2(n1663), .QN(n1617) );
  NAND2X0 U1684 ( .IN1(N171), .IN2(N511), .QN(n1663) );
  AND2X1 U1685 ( .IN1(n1664), .IN2(n1618), .Q(n1661) );
  NAND3X0 U1686 ( .IN1(n1665), .IN2(n1624), .IN3(n1666), .QN(n1618) );
  NAND2X0 U1687 ( .IN1(n1667), .IN2(n1668), .QN(n1666) );
  NAND3X0 U1688 ( .IN1(n1667), .IN2(n1668), .IN3(n1669), .QN(n1664) );
  NAND2X0 U1689 ( .IN1(n1665), .IN2(n1624), .QN(n1669) );
  AO21X1 U1690 ( .IN1(N188), .IN2(N494), .IN3(n1670), .Q(n1624) );
  NAND3X0 U1691 ( .IN1(N494), .IN2(n1670), .IN3(N188), .QN(n1665) );
  NAND2X0 U1692 ( .IN1(n1625), .IN2(n1671), .QN(n1670) );
  NAND3X0 U1693 ( .IN1(n1672), .IN2(n1673), .IN3(n1674), .QN(n1671) );
  AO21X1 U1694 ( .IN1(n1672), .IN2(n1673), .IN3(n1674), .Q(n1625) );
  NAND2X0 U1695 ( .IN1(n1630), .IN2(n1675), .QN(n1674) );
  NAND3X0 U1696 ( .IN1(N477), .IN2(n1676), .IN3(N205), .QN(n1675) );
  AO21X1 U1697 ( .IN1(N205), .IN2(N477), .IN3(n1676), .Q(n1630) );
  NAND2X0 U1698 ( .IN1(n1631), .IN2(n1677), .QN(n1676) );
  NAND3X0 U1699 ( .IN1(n1678), .IN2(n1679), .IN3(n1680), .QN(n1677) );
  AO21X1 U1700 ( .IN1(n1678), .IN2(n1679), .IN3(n1680), .Q(n1631) );
  NAND2X0 U1701 ( .IN1(n1637), .IN2(n1681), .QN(n1680) );
  NAND3X0 U1702 ( .IN1(N460), .IN2(n1682), .IN3(N222), .QN(n1681) );
  AO21X1 U1703 ( .IN1(N222), .IN2(N460), .IN3(n1682), .Q(n1637) );
  NAND2X0 U1704 ( .IN1(n1638), .IN2(n1683), .QN(n1682) );
  NAND3X0 U1705 ( .IN1(n1684), .IN2(n1685), .IN3(n1686), .QN(n1683) );
  AO21X1 U1706 ( .IN1(n1684), .IN2(n1685), .IN3(n1686), .Q(n1638) );
  NAND2X0 U1707 ( .IN1(n1603), .IN2(n1687), .QN(n1686) );
  NAND3X0 U1708 ( .IN1(N239), .IN2(n1688), .IN3(N443), .QN(n1687) );
  AO21X1 U1709 ( .IN1(N443), .IN2(N239), .IN3(n1688), .Q(n1603) );
  NAND2X0 U1710 ( .IN1(n1604), .IN2(n1689), .QN(n1688) );
  NAND3X0 U1711 ( .IN1(n1690), .IN2(n1691), .IN3(N426), .QN(n1689) );
  AO22X1 U1712 ( .IN1(N426), .IN2(N256), .IN3(n1690), .IN4(n1691), .Q(n1604)
         );
  NAND2X0 U1713 ( .IN1(n1645), .IN2(n1692), .QN(N6220) );
  NAND3X0 U1714 ( .IN1(n1693), .IN2(n1694), .IN3(n1695), .QN(n1692) );
  AO21X1 U1715 ( .IN1(n1693), .IN2(n1694), .IN3(n1695), .Q(n1645) );
  NAND2X0 U1716 ( .IN1(n1646), .IN2(n1696), .QN(n1695) );
  NAND3X0 U1717 ( .IN1(n1697), .IN2(n1698), .IN3(n1699), .QN(n1696) );
  AO21X1 U1718 ( .IN1(n1697), .IN2(n1698), .IN3(n1699), .Q(n1646) );
  NAND2X0 U1719 ( .IN1(n1649), .IN2(n1700), .QN(n1699) );
  NAND3X0 U1720 ( .IN1(N528), .IN2(n1701), .IN3(N137), .QN(n1700) );
  AO21X1 U1721 ( .IN1(N137), .IN2(N528), .IN3(n1701), .Q(n1649) );
  NAND2X0 U1722 ( .IN1(n1650), .IN2(n1702), .QN(n1701) );
  NAND3X0 U1723 ( .IN1(n1703), .IN2(n1704), .IN3(n1705), .QN(n1702) );
  AO21X1 U1724 ( .IN1(n1703), .IN2(n1704), .IN3(n1705), .Q(n1650) );
  NAND2X0 U1725 ( .IN1(n1660), .IN2(n1706), .QN(n1705) );
  NAND3X0 U1726 ( .IN1(N511), .IN2(n1707), .IN3(N154), .QN(n1706) );
  AO21X1 U1727 ( .IN1(N154), .IN2(N511), .IN3(n1707), .Q(n1660) );
  XNOR2X1 U1728 ( .IN1(n1658), .IN2(n1659), .Q(n1707) );
  AND2X1 U1729 ( .IN1(n1708), .IN2(n1709), .Q(n1659) );
  NAND2X0 U1730 ( .IN1(n1667), .IN2(n1710), .QN(n1658) );
  NAND3X0 U1731 ( .IN1(N494), .IN2(n1711), .IN3(N171), .QN(n1710) );
  AO21X1 U1732 ( .IN1(N171), .IN2(N494), .IN3(n1711), .Q(n1667) );
  NAND2X0 U1733 ( .IN1(n1668), .IN2(n1712), .QN(n1711) );
  NAND3X0 U1734 ( .IN1(n1713), .IN2(n1714), .IN3(n1715), .QN(n1712) );
  AO21X1 U1735 ( .IN1(n1713), .IN2(n1714), .IN3(n1715), .Q(n1668) );
  NAND2X0 U1736 ( .IN1(n1672), .IN2(n1716), .QN(n1715) );
  NAND3X0 U1737 ( .IN1(N477), .IN2(n1717), .IN3(N188), .QN(n1716) );
  AO21X1 U1738 ( .IN1(N188), .IN2(N477), .IN3(n1717), .Q(n1672) );
  NAND2X0 U1739 ( .IN1(n1673), .IN2(n1718), .QN(n1717) );
  NAND3X0 U1740 ( .IN1(n1719), .IN2(n1720), .IN3(n1721), .QN(n1718) );
  AO21X1 U1741 ( .IN1(n1719), .IN2(n1720), .IN3(n1721), .Q(n1673) );
  NAND2X0 U1742 ( .IN1(n1678), .IN2(n1722), .QN(n1721) );
  NAND3X0 U1743 ( .IN1(N460), .IN2(n1723), .IN3(N205), .QN(n1722) );
  AO21X1 U1744 ( .IN1(N205), .IN2(N460), .IN3(n1723), .Q(n1678) );
  NAND2X0 U1745 ( .IN1(n1679), .IN2(n1724), .QN(n1723) );
  NAND3X0 U1746 ( .IN1(n1725), .IN2(n1726), .IN3(n1727), .QN(n1724) );
  AO21X1 U1747 ( .IN1(n1725), .IN2(n1726), .IN3(n1727), .Q(n1679) );
  NAND2X0 U1748 ( .IN1(n1684), .IN2(n1728), .QN(n1727) );
  NAND3X0 U1749 ( .IN1(N443), .IN2(n1729), .IN3(N222), .QN(n1728) );
  AO21X1 U1750 ( .IN1(N222), .IN2(N443), .IN3(n1729), .Q(n1684) );
  NAND2X0 U1751 ( .IN1(n1685), .IN2(n1730), .QN(n1729) );
  NAND3X0 U1752 ( .IN1(n1731), .IN2(n1732), .IN3(n1733), .QN(n1730) );
  AO21X1 U1753 ( .IN1(n1731), .IN2(n1732), .IN3(n1733), .Q(n1685) );
  NAND2X0 U1754 ( .IN1(n1690), .IN2(n1734), .QN(n1733) );
  NAND3X0 U1755 ( .IN1(N239), .IN2(n1735), .IN3(N426), .QN(n1734) );
  AO21X1 U1756 ( .IN1(N426), .IN2(N239), .IN3(n1735), .Q(n1690) );
  AO21X1 U1757 ( .IN1(n1736), .IN2(N409), .IN3(n1737), .Q(n1735) );
  INVX0 U1758 ( .INP(n1691), .ZN(n1737) );
  AO21X1 U1759 ( .IN1(N409), .IN2(N256), .IN3(n1736), .Q(n1691) );
  AND2X1 U1760 ( .IN1(n1738), .IN2(n1739), .Q(n1736) );
  AO21X1 U1761 ( .IN1(N392), .IN2(N256), .IN3(n1740), .Q(n1738) );
  NAND2X0 U1762 ( .IN1(n1693), .IN2(n1741), .QN(N6210) );
  NAND3X0 U1763 ( .IN1(n1742), .IN2(n1743), .IN3(n1744), .QN(n1741) );
  AO21X1 U1764 ( .IN1(n1742), .IN2(n1743), .IN3(n1744), .Q(n1693) );
  AOI21X1 U1765 ( .IN1(n1694), .IN2(n1745), .IN3(n1746), .QN(n1744) );
  XOR2X1 U1766 ( .IN1(n1747), .IN2(keyinput29), .Q(n1746) );
  NAND2X0 U1767 ( .IN1(n1748), .IN2(n1694), .QN(n1747) );
  INVX0 U1768 ( .INP(n1749), .ZN(n1748) );
  NAND2X0 U1769 ( .IN1(n1750), .IN2(n1751), .QN(n1745) );
  AO21X1 U1770 ( .IN1(n1750), .IN2(n1751), .IN3(n1749), .Q(n1694) );
  NAND2X0 U1771 ( .IN1(n1697), .IN2(n1752), .QN(n1749) );
  NAND3X0 U1772 ( .IN1(N528), .IN2(n1753), .IN3(N120), .QN(n1752) );
  AO21X1 U1773 ( .IN1(N120), .IN2(N528), .IN3(n1753), .Q(n1697) );
  NAND2X0 U1774 ( .IN1(n1698), .IN2(n1754), .QN(n1753) );
  NAND3X0 U1775 ( .IN1(n1755), .IN2(n1756), .IN3(n1757), .QN(n1754) );
  AO21X1 U1776 ( .IN1(n1755), .IN2(n1756), .IN3(n1757), .Q(n1698) );
  NAND2X0 U1777 ( .IN1(n1703), .IN2(n1758), .QN(n1757) );
  NAND3X0 U1778 ( .IN1(N511), .IN2(n1759), .IN3(N137), .QN(n1758) );
  AO21X1 U1779 ( .IN1(N137), .IN2(N511), .IN3(n1759), .Q(n1703) );
  NAND2X0 U1780 ( .IN1(n1704), .IN2(n1760), .QN(n1759) );
  NAND3X0 U1781 ( .IN1(n1761), .IN2(n1762), .IN3(n1763), .QN(n1760) );
  AO21X1 U1782 ( .IN1(n1761), .IN2(n1762), .IN3(n1763), .Q(n1704) );
  NAND2X0 U1783 ( .IN1(n1709), .IN2(n1764), .QN(n1763) );
  NAND3X0 U1784 ( .IN1(N494), .IN2(n1765), .IN3(N154), .QN(n1764) );
  AO21X1 U1785 ( .IN1(N154), .IN2(N494), .IN3(n1765), .Q(n1709) );
  XNOR2X1 U1786 ( .IN1(n1766), .IN2(keyinput22), .Q(n1765) );
  NAND2X0 U1787 ( .IN1(n1708), .IN2(n1767), .QN(n1766) );
  NAND3X0 U1788 ( .IN1(n1768), .IN2(n1769), .IN3(n1770), .QN(n1767) );
  AO21X1 U1789 ( .IN1(n1768), .IN2(n1769), .IN3(n1770), .Q(n1708) );
  NAND2X0 U1790 ( .IN1(n1713), .IN2(n1771), .QN(n1770) );
  NAND3X0 U1791 ( .IN1(N477), .IN2(n1772), .IN3(N171), .QN(n1771) );
  AO21X1 U1792 ( .IN1(N171), .IN2(N477), .IN3(n1772), .Q(n1713) );
  NAND2X0 U1793 ( .IN1(n1714), .IN2(n1773), .QN(n1772) );
  NAND3X0 U1794 ( .IN1(n1774), .IN2(n1775), .IN3(n1776), .QN(n1773) );
  AO21X1 U1795 ( .IN1(n1774), .IN2(n1775), .IN3(n1776), .Q(n1714) );
  NAND2X0 U1796 ( .IN1(n1719), .IN2(n1777), .QN(n1776) );
  NAND3X0 U1797 ( .IN1(N460), .IN2(n1778), .IN3(N188), .QN(n1777) );
  AO21X1 U1798 ( .IN1(N188), .IN2(N460), .IN3(n1778), .Q(n1719) );
  NAND2X0 U1799 ( .IN1(n1720), .IN2(n1779), .QN(n1778) );
  NAND3X0 U1800 ( .IN1(n1780), .IN2(n1781), .IN3(n1782), .QN(n1779) );
  AO21X1 U1801 ( .IN1(n1780), .IN2(n1781), .IN3(n1782), .Q(n1720) );
  NAND2X0 U1802 ( .IN1(n1725), .IN2(n1783), .QN(n1782) );
  NAND3X0 U1803 ( .IN1(N443), .IN2(n1784), .IN3(N205), .QN(n1783) );
  AO21X1 U1804 ( .IN1(N205), .IN2(N443), .IN3(n1784), .Q(n1725) );
  NAND2X0 U1805 ( .IN1(n1726), .IN2(n1785), .QN(n1784) );
  NAND3X0 U1806 ( .IN1(n1786), .IN2(n1787), .IN3(n1788), .QN(n1785) );
  AO21X1 U1807 ( .IN1(n1786), .IN2(n1787), .IN3(n1788), .Q(n1726) );
  NAND2X0 U1808 ( .IN1(n1731), .IN2(n1789), .QN(n1788) );
  NAND3X0 U1809 ( .IN1(N426), .IN2(n1790), .IN3(N222), .QN(n1789) );
  AO21X1 U1810 ( .IN1(N222), .IN2(N426), .IN3(n1790), .Q(n1731) );
  NAND2X0 U1811 ( .IN1(n1732), .IN2(n1791), .QN(n1790) );
  NAND3X0 U1812 ( .IN1(n1792), .IN2(n1793), .IN3(n1794), .QN(n1791) );
  AO21X1 U1813 ( .IN1(n1792), .IN2(n1793), .IN3(n1794), .Q(n1732) );
  NAND2X0 U1814 ( .IN1(n1739), .IN2(n1795), .QN(n1794) );
  NAND3X0 U1815 ( .IN1(N409), .IN2(N239), .IN3(n1796), .QN(n1795) );
  AO21X1 U1816 ( .IN1(N409), .IN2(N239), .IN3(n1796), .Q(n1739) );
  XOR2X1 U1817 ( .IN1(n1797), .IN2(n1740), .Q(n1796) );
  AND2X1 U1818 ( .IN1(n1798), .IN2(n1799), .Q(n1740) );
  AO21X1 U1819 ( .IN1(N375), .IN2(N256), .IN3(n1800), .Q(n1798) );
  NAND2X0 U1820 ( .IN1(N392), .IN2(N256), .QN(n1797) );
  NAND2X0 U1821 ( .IN1(n1742), .IN2(n1801), .QN(N6200) );
  NAND3X0 U1822 ( .IN1(n1802), .IN2(n1803), .IN3(n1804), .QN(n1801) );
  AO21X1 U1823 ( .IN1(n1802), .IN2(n1803), .IN3(n1804), .Q(n1742) );
  NAND2X0 U1824 ( .IN1(n1743), .IN2(n1805), .QN(n1804) );
  NAND3X0 U1825 ( .IN1(n1806), .IN2(n1807), .IN3(n1808), .QN(n1805) );
  AO21X1 U1826 ( .IN1(n1806), .IN2(n1807), .IN3(n1808), .Q(n1743) );
  NAND2X0 U1827 ( .IN1(n1750), .IN2(n1809), .QN(n1808) );
  NAND3X0 U1828 ( .IN1(N528), .IN2(n1810), .IN3(N103), .QN(n1809) );
  AO21X1 U1829 ( .IN1(N103), .IN2(N528), .IN3(n1810), .Q(n1750) );
  NAND2X0 U1830 ( .IN1(n1751), .IN2(n1811), .QN(n1810) );
  NAND3X0 U1831 ( .IN1(n1812), .IN2(n1813), .IN3(n1814), .QN(n1811) );
  AO21X1 U1832 ( .IN1(n1812), .IN2(n1813), .IN3(n1814), .Q(n1751) );
  NAND2X0 U1833 ( .IN1(n1755), .IN2(n1815), .QN(n1814) );
  NAND3X0 U1834 ( .IN1(N511), .IN2(n1816), .IN3(N120), .QN(n1815) );
  AO21X1 U1835 ( .IN1(N120), .IN2(N511), .IN3(n1816), .Q(n1755) );
  NAND2X0 U1836 ( .IN1(n1756), .IN2(n1817), .QN(n1816) );
  NAND3X0 U1837 ( .IN1(n1818), .IN2(n1819), .IN3(n1820), .QN(n1817) );
  AO21X1 U1838 ( .IN1(n1818), .IN2(n1819), .IN3(n1820), .Q(n1756) );
  NAND2X0 U1839 ( .IN1(n1761), .IN2(n1821), .QN(n1820) );
  NAND3X0 U1840 ( .IN1(N137), .IN2(N494), .IN3(n1822), .QN(n1821) );
  AO21X1 U1841 ( .IN1(N137), .IN2(N494), .IN3(n1822), .Q(n1761) );
  AND2X1 U1842 ( .IN1(n1823), .IN2(n1824), .Q(n1822) );
  AO21X1 U1843 ( .IN1(n1825), .IN2(n1826), .IN3(n1827), .Q(n1824) );
  XOR2X1 U1844 ( .IN1(n1828), .IN2(keyinput21), .Q(n1823) );
  OR2X1 U1845 ( .IN1(n1829), .IN2(n1827), .Q(n1828) );
  INVX0 U1846 ( .INP(n1762), .ZN(n1827) );
  AO21X1 U1847 ( .IN1(n1825), .IN2(n1826), .IN3(n1829), .Q(n1762) );
  NAND2X0 U1848 ( .IN1(n1830), .IN2(n1768), .QN(n1829) );
  NAND3X0 U1849 ( .IN1(n1831), .IN2(n1769), .IN3(n1832), .QN(n1768) );
  NAND2X0 U1850 ( .IN1(N154), .IN2(N477), .QN(n1832) );
  NAND3X0 U1851 ( .IN1(N477), .IN2(n1833), .IN3(N154), .QN(n1830) );
  NAND2X0 U1852 ( .IN1(n1831), .IN2(n1769), .QN(n1833) );
  AO21X1 U1853 ( .IN1(n1834), .IN2(n1835), .IN3(n1836), .Q(n1769) );
  NAND3X0 U1854 ( .IN1(n1834), .IN2(n1835), .IN3(n1836), .QN(n1831) );
  NAND2X0 U1855 ( .IN1(n1774), .IN2(n1837), .QN(n1836) );
  NAND3X0 U1856 ( .IN1(N460), .IN2(n1838), .IN3(N171), .QN(n1837) );
  AO21X1 U1857 ( .IN1(N171), .IN2(N460), .IN3(n1838), .Q(n1774) );
  NAND2X0 U1858 ( .IN1(n1775), .IN2(n1839), .QN(n1838) );
  NAND3X0 U1859 ( .IN1(n1840), .IN2(n1841), .IN3(n1842), .QN(n1839) );
  AO21X1 U1860 ( .IN1(n1840), .IN2(n1841), .IN3(n1842), .Q(n1775) );
  NAND2X0 U1861 ( .IN1(n1780), .IN2(n1843), .QN(n1842) );
  NAND3X0 U1862 ( .IN1(N443), .IN2(n1844), .IN3(N188), .QN(n1843) );
  AO21X1 U1863 ( .IN1(N188), .IN2(N443), .IN3(n1844), .Q(n1780) );
  NAND2X0 U1864 ( .IN1(n1781), .IN2(n1845), .QN(n1844) );
  NAND3X0 U1865 ( .IN1(n1846), .IN2(n1847), .IN3(n1848), .QN(n1845) );
  AO21X1 U1866 ( .IN1(n1846), .IN2(n1847), .IN3(n1848), .Q(n1781) );
  NAND2X0 U1867 ( .IN1(n1786), .IN2(n1849), .QN(n1848) );
  NAND3X0 U1868 ( .IN1(N426), .IN2(n1850), .IN3(N205), .QN(n1849) );
  AO21X1 U1869 ( .IN1(N205), .IN2(N426), .IN3(n1850), .Q(n1786) );
  NAND2X0 U1870 ( .IN1(n1787), .IN2(n1851), .QN(n1850) );
  NAND3X0 U1871 ( .IN1(n1852), .IN2(n1853), .IN3(n1854), .QN(n1851) );
  AO21X1 U1872 ( .IN1(n1852), .IN2(n1853), .IN3(n1854), .Q(n1787) );
  NAND2X0 U1873 ( .IN1(n1792), .IN2(n1855), .QN(n1854) );
  NAND3X0 U1874 ( .IN1(N409), .IN2(n1856), .IN3(N222), .QN(n1855) );
  AO21X1 U1875 ( .IN1(N222), .IN2(N409), .IN3(n1856), .Q(n1792) );
  NAND2X0 U1876 ( .IN1(n1793), .IN2(n1857), .QN(n1856) );
  NAND3X0 U1877 ( .IN1(n1858), .IN2(n1859), .IN3(n1860), .QN(n1857) );
  AO21X1 U1878 ( .IN1(n1858), .IN2(n1859), .IN3(n1860), .Q(n1793) );
  NAND2X0 U1879 ( .IN1(n1799), .IN2(n1861), .QN(n1860) );
  NAND3X0 U1880 ( .IN1(N392), .IN2(N239), .IN3(n1862), .QN(n1861) );
  AO21X1 U1881 ( .IN1(N392), .IN2(N239), .IN3(n1862), .Q(n1799) );
  XOR2X1 U1882 ( .IN1(n1863), .IN2(n1800), .Q(n1862) );
  AND2X1 U1883 ( .IN1(n1864), .IN2(n1865), .Q(n1800) );
  AO21X1 U1884 ( .IN1(N358), .IN2(N256), .IN3(n1866), .Q(n1864) );
  NAND2X0 U1885 ( .IN1(N375), .IN2(N256), .QN(n1863) );
  NAND2X0 U1886 ( .IN1(n1802), .IN2(n1867), .QN(N6190) );
  NAND3X0 U1887 ( .IN1(n1868), .IN2(n1869), .IN3(n1870), .QN(n1867) );
  AO21X1 U1888 ( .IN1(n1868), .IN2(n1869), .IN3(n1870), .Q(n1802) );
  NAND2X0 U1889 ( .IN1(n1803), .IN2(n1871), .QN(n1870) );
  NAND3X0 U1890 ( .IN1(n1872), .IN2(n1873), .IN3(n1874), .QN(n1871) );
  AO21X1 U1891 ( .IN1(n1872), .IN2(n1873), .IN3(n1874), .Q(n1803) );
  NAND2X0 U1892 ( .IN1(n1806), .IN2(n1875), .QN(n1874) );
  NAND3X0 U1893 ( .IN1(N528), .IN2(n1876), .IN3(N86), .QN(n1875) );
  AO21X1 U1894 ( .IN1(N86), .IN2(N528), .IN3(n1876), .Q(n1806) );
  NAND2X0 U1895 ( .IN1(n1807), .IN2(n1877), .QN(n1876) );
  NAND3X0 U1896 ( .IN1(n1878), .IN2(n1879), .IN3(n1880), .QN(n1877) );
  AO21X1 U1897 ( .IN1(n1878), .IN2(n1879), .IN3(n1880), .Q(n1807) );
  NAND2X0 U1898 ( .IN1(n1812), .IN2(n1881), .QN(n1880) );
  NAND3X0 U1899 ( .IN1(N511), .IN2(n1882), .IN3(N103), .QN(n1881) );
  AO21X1 U1900 ( .IN1(N103), .IN2(N511), .IN3(n1882), .Q(n1812) );
  NAND2X0 U1901 ( .IN1(n1813), .IN2(n1883), .QN(n1882) );
  NAND3X0 U1902 ( .IN1(n1884), .IN2(n1885), .IN3(n1886), .QN(n1883) );
  AO21X1 U1903 ( .IN1(n1884), .IN2(n1885), .IN3(n1886), .Q(n1813) );
  NAND2X0 U1904 ( .IN1(n1818), .IN2(n1887), .QN(n1886) );
  NAND3X0 U1905 ( .IN1(N494), .IN2(n1888), .IN3(N120), .QN(n1887) );
  AO21X1 U1906 ( .IN1(N120), .IN2(N494), .IN3(n1888), .Q(n1818) );
  NAND2X0 U1907 ( .IN1(n1819), .IN2(n1889), .QN(n1888) );
  NAND3X0 U1908 ( .IN1(n1890), .IN2(n1891), .IN3(n1892), .QN(n1889) );
  AO21X1 U1909 ( .IN1(n1890), .IN2(n1891), .IN3(n1892), .Q(n1819) );
  NAND2X0 U1910 ( .IN1(n1825), .IN2(n1893), .QN(n1892) );
  NAND3X0 U1911 ( .IN1(N477), .IN2(n1894), .IN3(N137), .QN(n1893) );
  AO21X1 U1912 ( .IN1(N137), .IN2(N477), .IN3(n1894), .Q(n1825) );
  NAND2X0 U1913 ( .IN1(n1826), .IN2(n1895), .QN(n1894) );
  NAND3X0 U1914 ( .IN1(n1896), .IN2(n1897), .IN3(n1898), .QN(n1895) );
  AO21X1 U1915 ( .IN1(n1896), .IN2(n1897), .IN3(n1898), .Q(n1826) );
  NAND2X0 U1916 ( .IN1(n1834), .IN2(n1899), .QN(n1898) );
  NAND3X0 U1917 ( .IN1(N460), .IN2(n1900), .IN3(N154), .QN(n1899) );
  AO21X1 U1918 ( .IN1(N154), .IN2(N460), .IN3(n1900), .Q(n1834) );
  NAND2X0 U1919 ( .IN1(n1835), .IN2(n1901), .QN(n1900) );
  NAND3X0 U1920 ( .IN1(n1902), .IN2(n1903), .IN3(n1904), .QN(n1901) );
  AO21X1 U1921 ( .IN1(n1902), .IN2(n1903), .IN3(n1904), .Q(n1835) );
  NOR2X0 U1922 ( .IN1(n1905), .IN2(n1906), .QN(n1904) );
  INVX0 U1923 ( .INP(n1907), .ZN(n1906) );
  NAND2X0 U1924 ( .IN1(n1908), .IN2(n1840), .QN(n1903) );
  XNOR2X1 U1925 ( .IN1(n1909), .IN2(keyinput17), .Q(n1902) );
  NAND2X0 U1926 ( .IN1(n1840), .IN2(n1910), .QN(n1909) );
  NAND2X0 U1927 ( .IN1(n1908), .IN2(n1910), .QN(n1840) );
  NAND2X0 U1928 ( .IN1(N171), .IN2(N443), .QN(n1910) );
  AND2X1 U1929 ( .IN1(n1841), .IN2(n1911), .Q(n1908) );
  NAND3X0 U1930 ( .IN1(n1912), .IN2(n1913), .IN3(n1914), .QN(n1911) );
  AO21X1 U1931 ( .IN1(n1912), .IN2(n1913), .IN3(n1914), .Q(n1841) );
  NAND2X0 U1932 ( .IN1(n1846), .IN2(n1915), .QN(n1914) );
  NAND3X0 U1933 ( .IN1(N426), .IN2(n1916), .IN3(N188), .QN(n1915) );
  AO21X1 U1934 ( .IN1(N188), .IN2(N426), .IN3(n1916), .Q(n1846) );
  NAND2X0 U1935 ( .IN1(n1847), .IN2(n1917), .QN(n1916) );
  NAND3X0 U1936 ( .IN1(n1918), .IN2(n1919), .IN3(n1920), .QN(n1917) );
  AO21X1 U1937 ( .IN1(n1918), .IN2(n1919), .IN3(n1920), .Q(n1847) );
  NAND2X0 U1938 ( .IN1(n1852), .IN2(n1921), .QN(n1920) );
  NAND3X0 U1939 ( .IN1(N409), .IN2(n1922), .IN3(N205), .QN(n1921) );
  AO21X1 U1940 ( .IN1(N205), .IN2(N409), .IN3(n1922), .Q(n1852) );
  NAND2X0 U1941 ( .IN1(n1853), .IN2(n1923), .QN(n1922) );
  NAND3X0 U1942 ( .IN1(n1924), .IN2(n1925), .IN3(n1926), .QN(n1923) );
  AO21X1 U1943 ( .IN1(n1924), .IN2(n1925), .IN3(n1926), .Q(n1853) );
  NAND2X0 U1944 ( .IN1(n1858), .IN2(n1927), .QN(n1926) );
  NAND3X0 U1945 ( .IN1(N392), .IN2(n1928), .IN3(N222), .QN(n1927) );
  AO21X1 U1946 ( .IN1(N222), .IN2(N392), .IN3(n1928), .Q(n1858) );
  NAND2X0 U1947 ( .IN1(n1859), .IN2(n1929), .QN(n1928) );
  NAND3X0 U1948 ( .IN1(n1930), .IN2(n1931), .IN3(n1932), .QN(n1929) );
  AO21X1 U1949 ( .IN1(n1930), .IN2(n1931), .IN3(n1932), .Q(n1859) );
  AOI21X1 U1950 ( .IN1(n1933), .IN2(n1934), .IN3(n1935), .QN(n1932) );
  INVX0 U1951 ( .INP(n1936), .ZN(n1935) );
  NAND2X0 U1952 ( .IN1(n1937), .IN2(n1865), .QN(n1931) );
  XOR2X1 U1953 ( .IN1(n1938), .IN2(keyinput14), .Q(n1930) );
  NAND2X0 U1954 ( .IN1(n1865), .IN2(n1939), .QN(n1938) );
  NAND2X0 U1955 ( .IN1(n1937), .IN2(n1939), .QN(n1865) );
  NAND2X0 U1956 ( .IN1(N375), .IN2(N239), .QN(n1939) );
  XOR2X1 U1957 ( .IN1(n1866), .IN2(n1940), .Q(n1937) );
  AND2X1 U1958 ( .IN1(N256), .IN2(N358), .Q(n1940) );
  AND2X1 U1959 ( .IN1(n1941), .IN2(n1942), .Q(n1866) );
  AO21X1 U1960 ( .IN1(N341), .IN2(N256), .IN3(n1943), .Q(n1941) );
  NAND2X0 U1961 ( .IN1(n1868), .IN2(n1944), .QN(N6180) );
  NAND3X0 U1962 ( .IN1(n1945), .IN2(n1946), .IN3(n1947), .QN(n1944) );
  AO21X1 U1963 ( .IN1(n1945), .IN2(n1946), .IN3(n1947), .Q(n1868) );
  NAND2X0 U1964 ( .IN1(n1869), .IN2(n1948), .QN(n1947) );
  NAND3X0 U1965 ( .IN1(n1949), .IN2(n1950), .IN3(n1951), .QN(n1948) );
  AO21X1 U1966 ( .IN1(n1949), .IN2(n1950), .IN3(n1951), .Q(n1869) );
  NAND2X0 U1967 ( .IN1(n1872), .IN2(n1952), .QN(n1951) );
  NAND3X0 U1968 ( .IN1(N528), .IN2(n1953), .IN3(N69), .QN(n1952) );
  AO21X1 U1969 ( .IN1(N69), .IN2(N528), .IN3(n1953), .Q(n1872) );
  NAND2X0 U1970 ( .IN1(n1873), .IN2(n1954), .QN(n1953) );
  NAND3X0 U1971 ( .IN1(n1955), .IN2(n1956), .IN3(n1957), .QN(n1954) );
  AO21X1 U1972 ( .IN1(n1955), .IN2(n1956), .IN3(n1957), .Q(n1873) );
  NAND2X0 U1973 ( .IN1(n1878), .IN2(n1958), .QN(n1957) );
  NAND3X0 U1974 ( .IN1(N511), .IN2(n1959), .IN3(N86), .QN(n1958) );
  AO21X1 U1975 ( .IN1(N86), .IN2(N511), .IN3(n1959), .Q(n1878) );
  NAND2X0 U1976 ( .IN1(n1879), .IN2(n1960), .QN(n1959) );
  NAND4X0 U1977 ( .IN1(n1961), .IN2(n1962), .IN3(n1963), .IN4(n1964), .QN(
        n1960) );
  AO22X1 U1978 ( .IN1(n1963), .IN2(n1964), .IN3(n1961), .IN4(n1962), .Q(n1879)
         );
  AO21X1 U1979 ( .IN1(N103), .IN2(N494), .IN3(n1965), .Q(n1962) );
  XNOR2X1 U1980 ( .IN1(n1966), .IN2(keyinput23), .Q(n1961) );
  OR2X1 U1981 ( .IN1(n1967), .IN2(n1965), .Q(n1966) );
  INVX0 U1982 ( .INP(n1884), .ZN(n1965) );
  AO21X1 U1983 ( .IN1(N103), .IN2(N494), .IN3(n1967), .Q(n1884) );
  NAND2X0 U1984 ( .IN1(n1885), .IN2(n1968), .QN(n1967) );
  NAND3X0 U1985 ( .IN1(n1969), .IN2(n1970), .IN3(n1971), .QN(n1968) );
  AO21X1 U1986 ( .IN1(n1969), .IN2(n1970), .IN3(n1971), .Q(n1885) );
  NAND2X0 U1987 ( .IN1(n1890), .IN2(n1972), .QN(n1971) );
  NAND3X0 U1988 ( .IN1(N477), .IN2(n1973), .IN3(N120), .QN(n1972) );
  AO21X1 U1989 ( .IN1(N120), .IN2(N477), .IN3(n1973), .Q(n1890) );
  NAND2X0 U1990 ( .IN1(n1891), .IN2(n1974), .QN(n1973) );
  NAND3X0 U1991 ( .IN1(n1975), .IN2(n1976), .IN3(n1977), .QN(n1974) );
  AO21X1 U1992 ( .IN1(n1975), .IN2(n1976), .IN3(n1977), .Q(n1891) );
  NAND2X0 U1993 ( .IN1(n1896), .IN2(n1978), .QN(n1977) );
  NAND3X0 U1994 ( .IN1(N460), .IN2(n1979), .IN3(N137), .QN(n1978) );
  AO21X1 U1995 ( .IN1(N137), .IN2(N460), .IN3(n1979), .Q(n1896) );
  NAND2X0 U1996 ( .IN1(n1897), .IN2(n1980), .QN(n1979) );
  NAND3X0 U1997 ( .IN1(n1981), .IN2(n1982), .IN3(n1983), .QN(n1980) );
  AO21X1 U1998 ( .IN1(n1981), .IN2(n1982), .IN3(n1983), .Q(n1897) );
  AO21X1 U1999 ( .IN1(n1984), .IN2(n1985), .IN3(n1905), .Q(n1983) );
  NOR2X0 U2000 ( .IN1(n1985), .IN2(n1984), .QN(n1905) );
  NAND2X0 U2001 ( .IN1(n1907), .IN2(n1986), .QN(n1985) );
  NAND3X0 U2002 ( .IN1(n1987), .IN2(n1988), .IN3(n1989), .QN(n1986) );
  AO21X1 U2003 ( .IN1(n1987), .IN2(n1988), .IN3(n1989), .Q(n1907) );
  NAND2X0 U2004 ( .IN1(n1912), .IN2(n1990), .QN(n1989) );
  NAND3X0 U2005 ( .IN1(N426), .IN2(n1991), .IN3(N171), .QN(n1990) );
  AO21X1 U2006 ( .IN1(N171), .IN2(N426), .IN3(n1991), .Q(n1912) );
  NAND2X0 U2007 ( .IN1(n1913), .IN2(n1992), .QN(n1991) );
  NAND3X0 U2008 ( .IN1(n1993), .IN2(n1994), .IN3(n1995), .QN(n1992) );
  AO21X1 U2009 ( .IN1(n1993), .IN2(n1994), .IN3(n1995), .Q(n1913) );
  NAND2X0 U2010 ( .IN1(n1918), .IN2(n1996), .QN(n1995) );
  NAND3X0 U2011 ( .IN1(N409), .IN2(n1997), .IN3(N188), .QN(n1996) );
  AO21X1 U2012 ( .IN1(N188), .IN2(N409), .IN3(n1997), .Q(n1918) );
  NAND2X0 U2013 ( .IN1(n1919), .IN2(n1998), .QN(n1997) );
  NAND3X0 U2014 ( .IN1(n1999), .IN2(n2000), .IN3(n2001), .QN(n1998) );
  AO21X1 U2015 ( .IN1(n1999), .IN2(n2000), .IN3(n2001), .Q(n1919) );
  NAND2X0 U2016 ( .IN1(n1924), .IN2(n2002), .QN(n2001) );
  NAND3X0 U2017 ( .IN1(N392), .IN2(n2003), .IN3(N205), .QN(n2002) );
  AO21X1 U2018 ( .IN1(N205), .IN2(N392), .IN3(n2003), .Q(n1924) );
  NAND2X0 U2019 ( .IN1(n1925), .IN2(n2004), .QN(n2003) );
  NAND3X0 U2020 ( .IN1(n2005), .IN2(n2006), .IN3(n2007), .QN(n2004) );
  AO21X1 U2021 ( .IN1(n2005), .IN2(n2006), .IN3(n2007), .Q(n1925) );
  NAND2X0 U2022 ( .IN1(n1936), .IN2(n2008), .QN(n2007) );
  NAND3X0 U2023 ( .IN1(N375), .IN2(n2009), .IN3(N222), .QN(n2008) );
  AO21X1 U2024 ( .IN1(N222), .IN2(N375), .IN3(n2009), .Q(n1936) );
  XNOR2X1 U2025 ( .IN1(n1934), .IN2(n1933), .Q(n2009) );
  AND2X1 U2026 ( .IN1(n1942), .IN2(n2010), .Q(n1933) );
  NAND3X0 U2027 ( .IN1(N358), .IN2(N239), .IN3(n2011), .QN(n2010) );
  AO21X1 U2028 ( .IN1(N358), .IN2(N239), .IN3(n2011), .Q(n1942) );
  XNOR2X1 U2029 ( .IN1(n1943), .IN2(n2012), .Q(n2011) );
  AND2X1 U2030 ( .IN1(N256), .IN2(N341), .Q(n2012) );
  AOI21X1 U2031 ( .IN1(n2013), .IN2(n2014), .IN3(n2015), .QN(n1943) );
  INVX0 U2032 ( .INP(n2016), .ZN(n2015) );
  NAND2X0 U2033 ( .IN1(n2017), .IN2(n2018), .QN(n1934) );
  XNOR2X1 U2034 ( .IN1(n2019), .IN2(keyinput1), .Q(n1984) );
  NAND2X0 U2035 ( .IN1(N154), .IN2(N443), .QN(n2019) );
  NAND2X0 U2036 ( .IN1(n1945), .IN2(n2020), .QN(N6170) );
  AO221X1 U2037 ( .IN1(n2021), .IN2(n1946), .IN3(n2022), .IN4(n2023), .IN5(
        n2024), .Q(n2020) );
  NAND3X0 U2038 ( .IN1(n2021), .IN2(n1946), .IN3(n2025), .QN(n1945) );
  AO21X1 U2039 ( .IN1(n2022), .IN2(n2023), .IN3(n2024), .Q(n2025) );
  INVX0 U2040 ( .INP(n2026), .ZN(n2024) );
  AO21X1 U2041 ( .IN1(n2027), .IN2(n2028), .IN3(n2029), .Q(n1946) );
  NAND3X0 U2042 ( .IN1(n2027), .IN2(n2028), .IN3(n2029), .QN(n2021) );
  NAND2X0 U2043 ( .IN1(n1949), .IN2(n2030), .QN(n2029) );
  NAND3X0 U2044 ( .IN1(N528), .IN2(n2031), .IN3(N52), .QN(n2030) );
  AO21X1 U2045 ( .IN1(N52), .IN2(N528), .IN3(n2031), .Q(n1949) );
  NAND2X0 U2046 ( .IN1(n1950), .IN2(n2032), .QN(n2031) );
  NAND3X0 U2047 ( .IN1(n2033), .IN2(n2034), .IN3(n2035), .QN(n2032) );
  AO21X1 U2048 ( .IN1(n2033), .IN2(n2034), .IN3(n2035), .Q(n1950) );
  NAND2X0 U2049 ( .IN1(n1955), .IN2(n2036), .QN(n2035) );
  NAND3X0 U2050 ( .IN1(N511), .IN2(n2037), .IN3(N69), .QN(n2036) );
  AO21X1 U2051 ( .IN1(N69), .IN2(N511), .IN3(n2037), .Q(n1955) );
  NAND2X0 U2052 ( .IN1(n1956), .IN2(n2038), .QN(n2037) );
  NAND3X0 U2053 ( .IN1(n2039), .IN2(n2040), .IN3(n2041), .QN(n2038) );
  AO21X1 U2054 ( .IN1(n2039), .IN2(n2040), .IN3(n2041), .Q(n1956) );
  NAND2X0 U2055 ( .IN1(n1963), .IN2(n2042), .QN(n2041) );
  NAND3X0 U2056 ( .IN1(N494), .IN2(n2043), .IN3(N86), .QN(n2042) );
  AO21X1 U2057 ( .IN1(N86), .IN2(N494), .IN3(n2043), .Q(n1963) );
  NAND2X0 U2058 ( .IN1(n1964), .IN2(n2044), .QN(n2043) );
  NAND3X0 U2059 ( .IN1(n2045), .IN2(n2046), .IN3(n2047), .QN(n2044) );
  AO21X1 U2060 ( .IN1(n2045), .IN2(n2046), .IN3(n2047), .Q(n1964) );
  NAND2X0 U2061 ( .IN1(n1969), .IN2(n2048), .QN(n2047) );
  NAND3X0 U2062 ( .IN1(N477), .IN2(n2049), .IN3(N103), .QN(n2048) );
  AO21X1 U2063 ( .IN1(N103), .IN2(N477), .IN3(n2049), .Q(n1969) );
  NAND2X0 U2064 ( .IN1(n1970), .IN2(n2050), .QN(n2049) );
  NAND3X0 U2065 ( .IN1(n2051), .IN2(n2052), .IN3(n2053), .QN(n2050) );
  AO21X1 U2066 ( .IN1(n2051), .IN2(n2052), .IN3(n2053), .Q(n1970) );
  NAND2X0 U2067 ( .IN1(n1975), .IN2(n2054), .QN(n2053) );
  NAND3X0 U2068 ( .IN1(N460), .IN2(n2055), .IN3(N120), .QN(n2054) );
  AO21X1 U2069 ( .IN1(N120), .IN2(N460), .IN3(n2055), .Q(n1975) );
  NAND2X0 U2070 ( .IN1(n1976), .IN2(n2056), .QN(n2055) );
  NAND3X0 U2071 ( .IN1(n2057), .IN2(n2058), .IN3(n2059), .QN(n2056) );
  AO21X1 U2072 ( .IN1(n2057), .IN2(n2058), .IN3(n2059), .Q(n1976) );
  NAND2X0 U2073 ( .IN1(n1981), .IN2(n2060), .QN(n2059) );
  NAND3X0 U2074 ( .IN1(N443), .IN2(n2061), .IN3(N137), .QN(n2060) );
  AO21X1 U2075 ( .IN1(N137), .IN2(N443), .IN3(n2061), .Q(n1981) );
  NAND2X0 U2076 ( .IN1(n1982), .IN2(n2062), .QN(n2061) );
  NAND3X0 U2077 ( .IN1(n2063), .IN2(n2064), .IN3(n2065), .QN(n2062) );
  AO21X1 U2078 ( .IN1(n2063), .IN2(n2064), .IN3(n2065), .Q(n1982) );
  NAND2X0 U2079 ( .IN1(n1987), .IN2(n2066), .QN(n2065) );
  NAND3X0 U2080 ( .IN1(N426), .IN2(n2067), .IN3(N154), .QN(n2066) );
  AO21X1 U2081 ( .IN1(N154), .IN2(N426), .IN3(n2067), .Q(n1987) );
  NAND2X0 U2082 ( .IN1(n1988), .IN2(n2068), .QN(n2067) );
  NAND3X0 U2083 ( .IN1(n2069), .IN2(n2070), .IN3(n2071), .QN(n2068) );
  AO21X1 U2084 ( .IN1(n2069), .IN2(n2070), .IN3(n2071), .Q(n1988) );
  NAND2X0 U2085 ( .IN1(n1993), .IN2(n2072), .QN(n2071) );
  NAND3X0 U2086 ( .IN1(N409), .IN2(n2073), .IN3(N171), .QN(n2072) );
  AO21X1 U2087 ( .IN1(N171), .IN2(N409), .IN3(n2073), .Q(n1993) );
  NAND2X0 U2088 ( .IN1(n1994), .IN2(n2074), .QN(n2073) );
  NAND3X0 U2089 ( .IN1(n2075), .IN2(n2076), .IN3(n2077), .QN(n2074) );
  AO21X1 U2090 ( .IN1(n2075), .IN2(n2076), .IN3(n2077), .Q(n1994) );
  NAND2X0 U2091 ( .IN1(n1999), .IN2(n2078), .QN(n2077) );
  NAND3X0 U2092 ( .IN1(N392), .IN2(n2079), .IN3(N188), .QN(n2078) );
  AO21X1 U2093 ( .IN1(N188), .IN2(N392), .IN3(n2079), .Q(n1999) );
  NAND2X0 U2094 ( .IN1(n2000), .IN2(n2080), .QN(n2079) );
  NAND3X0 U2095 ( .IN1(n2081), .IN2(n2082), .IN3(n2083), .QN(n2080) );
  AO21X1 U2096 ( .IN1(n2081), .IN2(n2082), .IN3(n2083), .Q(n2000) );
  NAND2X0 U2097 ( .IN1(n2005), .IN2(n2084), .QN(n2083) );
  NAND4X0 U2098 ( .IN1(N205), .IN2(N375), .IN3(n2085), .IN4(n2086), .QN(n2084)
         );
  AO22X1 U2099 ( .IN1(N205), .IN2(N375), .IN3(n2085), .IN4(n2086), .Q(n2005)
         );
  OR2X1 U2100 ( .IN1(n2087), .IN2(n2088), .Q(n2086) );
  XOR2X1 U2101 ( .IN1(keyinput13), .IN2(n2089), .Q(n2085) );
  AOI21X1 U2102 ( .IN1(n2090), .IN2(n2091), .IN3(n2088), .QN(n2089) );
  INVX0 U2103 ( .INP(n2006), .ZN(n2088) );
  AO21X1 U2104 ( .IN1(n2091), .IN2(n2090), .IN3(n2087), .Q(n2006) );
  NAND2X0 U2105 ( .IN1(n2018), .IN2(n2092), .QN(n2087) );
  NAND3X0 U2106 ( .IN1(N358), .IN2(n2093), .IN3(N222), .QN(n2092) );
  AO21X1 U2107 ( .IN1(N222), .IN2(N358), .IN3(n2093), .Q(n2018) );
  NAND2X0 U2108 ( .IN1(n2017), .IN2(n2094), .QN(n2093) );
  NAND3X0 U2109 ( .IN1(n2095), .IN2(n2096), .IN3(n2097), .QN(n2094) );
  AO21X1 U2110 ( .IN1(n2095), .IN2(n2096), .IN3(n2097), .Q(n2017) );
  NAND2X0 U2111 ( .IN1(n2016), .IN2(n2098), .QN(n2097) );
  NAND3X0 U2112 ( .IN1(N341), .IN2(N239), .IN3(n2099), .QN(n2098) );
  AO21X1 U2113 ( .IN1(N341), .IN2(N239), .IN3(n2099), .Q(n2016) );
  XNOR2X1 U2114 ( .IN1(n2013), .IN2(n2014), .Q(n2099) );
  AO21X1 U2115 ( .IN1(n2100), .IN2(n2101), .IN3(n2102), .Q(n2014) );
  NAND2X0 U2116 ( .IN1(N324), .IN2(N256), .QN(n2013) );
  XNOR2X1 U2117 ( .IN1(n2023), .IN2(n2022), .Q(N6160) );
  AND2X1 U2118 ( .IN1(n2026), .IN2(n2103), .Q(n2022) );
  NAND3X0 U2119 ( .IN1(n2104), .IN2(n2105), .IN3(n2106), .QN(n2103) );
  AO21X1 U2120 ( .IN1(n2106), .IN2(n2104), .IN3(n2105), .Q(n2026) );
  NAND2X0 U2121 ( .IN1(n2027), .IN2(n2107), .QN(n2105) );
  NAND3X0 U2122 ( .IN1(N528), .IN2(n2108), .IN3(N35), .QN(n2107) );
  AO21X1 U2123 ( .IN1(N35), .IN2(N528), .IN3(n2108), .Q(n2027) );
  NAND2X0 U2124 ( .IN1(n2028), .IN2(n2109), .QN(n2108) );
  NAND3X0 U2125 ( .IN1(n2110), .IN2(n2111), .IN3(n2112), .QN(n2109) );
  AO21X1 U2126 ( .IN1(n2112), .IN2(n2111), .IN3(n2110), .Q(n2028) );
  NAND2X0 U2127 ( .IN1(n2033), .IN2(n2113), .QN(n2110) );
  NAND3X0 U2128 ( .IN1(N511), .IN2(n2114), .IN3(N52), .QN(n2113) );
  AO21X1 U2129 ( .IN1(N52), .IN2(N511), .IN3(n2114), .Q(n2033) );
  NAND2X0 U2130 ( .IN1(n2034), .IN2(n2115), .QN(n2114) );
  NAND3X0 U2131 ( .IN1(n2116), .IN2(n2117), .IN3(n2118), .QN(n2115) );
  AO21X1 U2132 ( .IN1(n2116), .IN2(n2117), .IN3(n2118), .Q(n2034) );
  NAND2X0 U2133 ( .IN1(n2039), .IN2(n2119), .QN(n2118) );
  NAND3X0 U2134 ( .IN1(N494), .IN2(n2120), .IN3(N69), .QN(n2119) );
  AO21X1 U2135 ( .IN1(N69), .IN2(N494), .IN3(n2120), .Q(n2039) );
  NAND2X0 U2136 ( .IN1(n2040), .IN2(n2121), .QN(n2120) );
  NAND3X0 U2137 ( .IN1(n2122), .IN2(n2123), .IN3(n2124), .QN(n2121) );
  AO21X1 U2138 ( .IN1(n2122), .IN2(n2123), .IN3(n2124), .Q(n2040) );
  NAND2X0 U2139 ( .IN1(n2045), .IN2(n2125), .QN(n2124) );
  NAND3X0 U2140 ( .IN1(N477), .IN2(n2126), .IN3(N86), .QN(n2125) );
  AO21X1 U2141 ( .IN1(N86), .IN2(N477), .IN3(n2126), .Q(n2045) );
  NAND2X0 U2142 ( .IN1(n2046), .IN2(n2127), .QN(n2126) );
  NAND3X0 U2143 ( .IN1(n2128), .IN2(n2129), .IN3(n2130), .QN(n2127) );
  AO21X1 U2144 ( .IN1(n2128), .IN2(n2129), .IN3(n2130), .Q(n2046) );
  NAND2X0 U2145 ( .IN1(n2051), .IN2(n2131), .QN(n2130) );
  NAND3X0 U2146 ( .IN1(N460), .IN2(n2132), .IN3(N103), .QN(n2131) );
  AO21X1 U2147 ( .IN1(N103), .IN2(N460), .IN3(n2132), .Q(n2051) );
  NAND2X0 U2148 ( .IN1(n2052), .IN2(n2133), .QN(n2132) );
  NAND3X0 U2149 ( .IN1(n2134), .IN2(n2135), .IN3(n2136), .QN(n2133) );
  AO21X1 U2150 ( .IN1(n2134), .IN2(n2135), .IN3(n2136), .Q(n2052) );
  NAND2X0 U2151 ( .IN1(n2057), .IN2(n2137), .QN(n2136) );
  NAND3X0 U2152 ( .IN1(N443), .IN2(n2138), .IN3(N120), .QN(n2137) );
  AO21X1 U2153 ( .IN1(N120), .IN2(N443), .IN3(n2138), .Q(n2057) );
  NAND2X0 U2154 ( .IN1(n2058), .IN2(n2139), .QN(n2138) );
  NAND3X0 U2155 ( .IN1(n2140), .IN2(n2141), .IN3(n2142), .QN(n2139) );
  AO21X1 U2156 ( .IN1(n2140), .IN2(n2141), .IN3(n2142), .Q(n2058) );
  NAND2X0 U2157 ( .IN1(n2063), .IN2(n2143), .QN(n2142) );
  NAND3X0 U2158 ( .IN1(N426), .IN2(n2144), .IN3(N137), .QN(n2143) );
  AO21X1 U2159 ( .IN1(N137), .IN2(N426), .IN3(n2144), .Q(n2063) );
  NAND2X0 U2160 ( .IN1(n2064), .IN2(n2145), .QN(n2144) );
  NAND3X0 U2161 ( .IN1(n2146), .IN2(n2147), .IN3(n2148), .QN(n2145) );
  AO21X1 U2162 ( .IN1(n2146), .IN2(n2147), .IN3(n2148), .Q(n2064) );
  NAND2X0 U2163 ( .IN1(n2069), .IN2(n2149), .QN(n2148) );
  NAND3X0 U2164 ( .IN1(N409), .IN2(n2150), .IN3(N154), .QN(n2149) );
  AO21X1 U2165 ( .IN1(N154), .IN2(N409), .IN3(n2150), .Q(n2069) );
  NAND2X0 U2166 ( .IN1(n2070), .IN2(n2151), .QN(n2150) );
  NAND3X0 U2167 ( .IN1(n2152), .IN2(n2153), .IN3(n2154), .QN(n2151) );
  AO21X1 U2168 ( .IN1(n2152), .IN2(n2153), .IN3(n2154), .Q(n2070) );
  NAND2X0 U2169 ( .IN1(n2075), .IN2(n2155), .QN(n2154) );
  NAND3X0 U2170 ( .IN1(N392), .IN2(n2156), .IN3(N171), .QN(n2155) );
  AO21X1 U2171 ( .IN1(N171), .IN2(N392), .IN3(n2156), .Q(n2075) );
  NAND2X0 U2172 ( .IN1(n2076), .IN2(n2157), .QN(n2156) );
  NAND3X0 U2173 ( .IN1(n2158), .IN2(n2159), .IN3(n2160), .QN(n2157) );
  AO21X1 U2174 ( .IN1(n2158), .IN2(n2159), .IN3(n2160), .Q(n2076) );
  NAND2X0 U2175 ( .IN1(n2081), .IN2(n2161), .QN(n2160) );
  NAND3X0 U2176 ( .IN1(N375), .IN2(n2162), .IN3(N188), .QN(n2161) );
  AO21X1 U2177 ( .IN1(N188), .IN2(N375), .IN3(n2162), .Q(n2081) );
  NAND2X0 U2178 ( .IN1(n2082), .IN2(n2163), .QN(n2162) );
  NAND3X0 U2179 ( .IN1(n2164), .IN2(n2165), .IN3(n2166), .QN(n2163) );
  AO21X1 U2180 ( .IN1(n2164), .IN2(n2165), .IN3(n2166), .Q(n2082) );
  NAND2X0 U2181 ( .IN1(n2091), .IN2(n2167), .QN(n2166) );
  NAND3X0 U2182 ( .IN1(N358), .IN2(n2168), .IN3(N205), .QN(n2167) );
  AO21X1 U2183 ( .IN1(N205), .IN2(N358), .IN3(n2168), .Q(n2091) );
  NAND2X0 U2184 ( .IN1(n2090), .IN2(n2169), .QN(n2168) );
  NAND3X0 U2185 ( .IN1(n2170), .IN2(n2171), .IN3(n2172), .QN(n2169) );
  AO21X1 U2186 ( .IN1(n2170), .IN2(n2171), .IN3(n2172), .Q(n2090) );
  NAND2X0 U2187 ( .IN1(n2095), .IN2(n2173), .QN(n2172) );
  NAND3X0 U2188 ( .IN1(N341), .IN2(n2174), .IN3(N222), .QN(n2173) );
  AO21X1 U2189 ( .IN1(N222), .IN2(N341), .IN3(n2174), .Q(n2095) );
  NAND2X0 U2190 ( .IN1(n2096), .IN2(n2175), .QN(n2174) );
  NAND3X0 U2191 ( .IN1(n2176), .IN2(n2177), .IN3(n2178), .QN(n2175) );
  AO21X1 U2192 ( .IN1(n2176), .IN2(n2177), .IN3(n2178), .Q(n2096) );
  XNOR2X1 U2193 ( .IN1(n2100), .IN2(n2101), .Q(n2178) );
  AO21X1 U2194 ( .IN1(n2179), .IN2(n2180), .IN3(n2181), .Q(n2101) );
  XOR2X1 U2195 ( .IN1(n2182), .IN2(keyinput8), .Q(n2181) );
  NAND2X0 U2196 ( .IN1(n2183), .IN2(n2179), .QN(n2182) );
  INVX0 U2197 ( .INP(n2102), .ZN(n2179) );
  OA21X1 U2198 ( .IN1(n2180), .IN2(n1502), .IN3(n2183), .Q(n2102) );
  INVX0 U2199 ( .INP(N256), .ZN(n1502) );
  INVX0 U2200 ( .INP(N307), .ZN(n2180) );
  NAND2X0 U2201 ( .IN1(N324), .IN2(N239), .QN(n2100) );
  INVX0 U2202 ( .INP(n2184), .ZN(n2106) );
  NOR2X0 U2203 ( .IN1(n2185), .IN2(n2186), .QN(N6150) );
  AOI221X1 U2204 ( .IN1(n2187), .IN2(n2188), .IN3(n2189), .IN4(n2190), .IN5(
        n2184), .QN(n2186) );
  INVX0 U2205 ( .INP(n2023), .ZN(n2185) );
  NAND3X0 U2206 ( .IN1(n2188), .IN2(n2187), .IN3(n2191), .QN(n2023) );
  AO21X1 U2207 ( .IN1(n2190), .IN2(n2189), .IN3(n2184), .Q(n2191) );
  XNOR2X1 U2208 ( .IN1(n2192), .IN2(keyinput31), .Q(n2184) );
  OR2X1 U2209 ( .IN1(n2189), .IN2(n2190), .Q(n2192) );
  NAND2X0 U2210 ( .IN1(n2104), .IN2(n2193), .QN(n2189) );
  NAND3X0 U2211 ( .IN1(n2194), .IN2(n2195), .IN3(n2196), .QN(n2193) );
  XOR2X1 U2212 ( .IN1(keyinput28), .IN2(n2197), .Q(n2104) );
  AOI21X1 U2213 ( .IN1(n2194), .IN2(n2196), .IN3(n2195), .QN(n2197) );
  OAI21X1 U2214 ( .IN1(n2198), .IN2(n2199), .IN3(n2112), .QN(n2195) );
  XNOR2X1 U2215 ( .IN1(n2200), .IN2(keyinput27), .Q(n2112) );
  NAND2X0 U2216 ( .IN1(n2199), .IN2(n2198), .QN(n2200) );
  AND2X1 U2217 ( .IN1(n2111), .IN2(n2201), .Q(n2199) );
  NAND3X0 U2218 ( .IN1(n2202), .IN2(n2203), .IN3(n2204), .QN(n2201) );
  AO21X1 U2219 ( .IN1(n2202), .IN2(n2203), .IN3(n2204), .Q(n2111) );
  NAND2X0 U2220 ( .IN1(n2116), .IN2(n2205), .QN(n2204) );
  NAND3X0 U2221 ( .IN1(N494), .IN2(n2206), .IN3(N52), .QN(n2205) );
  AO21X1 U2222 ( .IN1(N52), .IN2(N494), .IN3(n2206), .Q(n2116) );
  NAND2X0 U2223 ( .IN1(n2117), .IN2(n2207), .QN(n2206) );
  NAND3X0 U2224 ( .IN1(n2208), .IN2(n2209), .IN3(n2210), .QN(n2207) );
  AO21X1 U2225 ( .IN1(n2208), .IN2(n2209), .IN3(n2210), .Q(n2117) );
  NAND2X0 U2226 ( .IN1(n2122), .IN2(n2211), .QN(n2210) );
  NAND3X0 U2227 ( .IN1(N477), .IN2(n2212), .IN3(N69), .QN(n2211) );
  AO21X1 U2228 ( .IN1(N69), .IN2(N477), .IN3(n2212), .Q(n2122) );
  NAND2X0 U2229 ( .IN1(n2123), .IN2(n2213), .QN(n2212) );
  NAND3X0 U2230 ( .IN1(n2214), .IN2(n2215), .IN3(n2216), .QN(n2213) );
  AO21X1 U2231 ( .IN1(n2216), .IN2(n2215), .IN3(n2214), .Q(n2123) );
  NAND2X0 U2232 ( .IN1(n2128), .IN2(n2217), .QN(n2214) );
  NAND3X0 U2233 ( .IN1(N460), .IN2(n2218), .IN3(N86), .QN(n2217) );
  AO21X1 U2234 ( .IN1(N86), .IN2(N460), .IN3(n2218), .Q(n2128) );
  NAND2X0 U2235 ( .IN1(n2129), .IN2(n2219), .QN(n2218) );
  NAND3X0 U2236 ( .IN1(n2220), .IN2(n2221), .IN3(n2222), .QN(n2219) );
  AO21X1 U2237 ( .IN1(n2220), .IN2(n2221), .IN3(n2222), .Q(n2129) );
  NAND2X0 U2238 ( .IN1(n2134), .IN2(n2223), .QN(n2222) );
  NAND3X0 U2239 ( .IN1(N443), .IN2(n2224), .IN3(N103), .QN(n2223) );
  AO21X1 U2240 ( .IN1(N103), .IN2(N443), .IN3(n2224), .Q(n2134) );
  NAND2X0 U2241 ( .IN1(n2135), .IN2(n2225), .QN(n2224) );
  NAND3X0 U2242 ( .IN1(n2226), .IN2(n2227), .IN3(n2228), .QN(n2225) );
  AO21X1 U2243 ( .IN1(n2226), .IN2(n2227), .IN3(n2228), .Q(n2135) );
  NAND2X0 U2244 ( .IN1(n2140), .IN2(n2229), .QN(n2228) );
  NAND3X0 U2245 ( .IN1(N426), .IN2(n2230), .IN3(N120), .QN(n2229) );
  AO21X1 U2246 ( .IN1(N120), .IN2(N426), .IN3(n2230), .Q(n2140) );
  NAND2X0 U2247 ( .IN1(n2141), .IN2(n2231), .QN(n2230) );
  NAND3X0 U2248 ( .IN1(n2232), .IN2(n2233), .IN3(n2234), .QN(n2231) );
  AO21X1 U2249 ( .IN1(n2232), .IN2(n2233), .IN3(n2234), .Q(n2141) );
  NAND2X0 U2250 ( .IN1(n2146), .IN2(n2235), .QN(n2234) );
  NAND3X0 U2251 ( .IN1(N409), .IN2(n2236), .IN3(N137), .QN(n2235) );
  AO21X1 U2252 ( .IN1(N137), .IN2(N409), .IN3(n2236), .Q(n2146) );
  NAND2X0 U2253 ( .IN1(n2147), .IN2(n2237), .QN(n2236) );
  NAND3X0 U2254 ( .IN1(n2238), .IN2(n2239), .IN3(n2240), .QN(n2237) );
  AO21X1 U2255 ( .IN1(n2238), .IN2(n2239), .IN3(n2240), .Q(n2147) );
  NAND2X0 U2256 ( .IN1(n2152), .IN2(n2241), .QN(n2240) );
  NAND3X0 U2257 ( .IN1(N392), .IN2(n2242), .IN3(N154), .QN(n2241) );
  AO21X1 U2258 ( .IN1(N154), .IN2(N392), .IN3(n2242), .Q(n2152) );
  NAND2X0 U2259 ( .IN1(n2153), .IN2(n2243), .QN(n2242) );
  NAND3X0 U2260 ( .IN1(n2244), .IN2(n2245), .IN3(n2246), .QN(n2243) );
  AO21X1 U2261 ( .IN1(n2244), .IN2(n2245), .IN3(n2246), .Q(n2153) );
  NAND2X0 U2262 ( .IN1(n2158), .IN2(n2247), .QN(n2246) );
  NAND3X0 U2263 ( .IN1(N375), .IN2(n2248), .IN3(N171), .QN(n2247) );
  AO21X1 U2264 ( .IN1(N171), .IN2(N375), .IN3(n2248), .Q(n2158) );
  NAND2X0 U2265 ( .IN1(n2159), .IN2(n2249), .QN(n2248) );
  NAND3X0 U2266 ( .IN1(n2250), .IN2(n2251), .IN3(n2252), .QN(n2249) );
  AO21X1 U2267 ( .IN1(n2250), .IN2(n2251), .IN3(n2252), .Q(n2159) );
  NAND2X0 U2268 ( .IN1(n2164), .IN2(n2253), .QN(n2252) );
  NAND3X0 U2269 ( .IN1(N358), .IN2(n2254), .IN3(N188), .QN(n2253) );
  AO21X1 U2270 ( .IN1(N188), .IN2(N358), .IN3(n2254), .Q(n2164) );
  NAND2X0 U2271 ( .IN1(n2165), .IN2(n2255), .QN(n2254) );
  NAND3X0 U2272 ( .IN1(n2256), .IN2(n2257), .IN3(n2258), .QN(n2255) );
  AO21X1 U2273 ( .IN1(n2256), .IN2(n2257), .IN3(n2258), .Q(n2165) );
  NAND2X0 U2274 ( .IN1(n2170), .IN2(n2259), .QN(n2258) );
  NAND3X0 U2275 ( .IN1(N341), .IN2(n2260), .IN3(N205), .QN(n2259) );
  AO21X1 U2276 ( .IN1(N205), .IN2(N341), .IN3(n2260), .Q(n2170) );
  NAND2X0 U2277 ( .IN1(n2171), .IN2(n2261), .QN(n2260) );
  NAND3X0 U2278 ( .IN1(n2262), .IN2(n2263), .IN3(n2264), .QN(n2261) );
  AO21X1 U2279 ( .IN1(n2262), .IN2(n2263), .IN3(n2264), .Q(n2171) );
  NAND2X0 U2280 ( .IN1(n2176), .IN2(n2265), .QN(n2264) );
  NAND3X0 U2281 ( .IN1(N324), .IN2(n2266), .IN3(N222), .QN(n2265) );
  AO21X1 U2282 ( .IN1(N222), .IN2(N324), .IN3(n2266), .Q(n2176) );
  NAND2X0 U2283 ( .IN1(n2177), .IN2(n2267), .QN(n2266) );
  NAND3X0 U2284 ( .IN1(n2268), .IN2(n2269), .IN3(n2270), .QN(n2267) );
  AO21X1 U2285 ( .IN1(n2268), .IN2(n2269), .IN3(n2270), .Q(n2177) );
  AND2X1 U2286 ( .IN1(n2271), .IN2(n2272), .Q(n2270) );
  NAND2X0 U2287 ( .IN1(n2273), .IN2(n2274), .QN(n2269) );
  INVX0 U2288 ( .INP(n2183), .ZN(n2273) );
  NAND3X0 U2289 ( .IN1(N256), .IN2(n2275), .IN3(N290), .QN(n2183) );
  XOR2X1 U2290 ( .IN1(n2276), .IN2(keyinput7), .Q(n2268) );
  NAND2X0 U2291 ( .IN1(n2275), .IN2(n2277), .QN(n2276) );
  NAND4X0 U2292 ( .IN1(N290), .IN2(N256), .IN3(n2277), .IN4(n2274), .QN(n2275)
         );
  NAND2X0 U2293 ( .IN1(N307), .IN2(N239), .QN(n2277) );
  NAND2X0 U2294 ( .IN1(N35), .IN2(N511), .QN(n2198) );
  AND2X1 U2295 ( .IN1(N18), .IN2(N528), .Q(n2190) );
  NAND2X0 U2296 ( .IN1(n2188), .IN2(n2278), .QN(N6123) );
  NAND3X0 U2297 ( .IN1(N528), .IN2(n2279), .IN3(N1), .QN(n2278) );
  AO21X1 U2298 ( .IN1(N1), .IN2(N528), .IN3(n2279), .Q(n2188) );
  XNOR2X1 U2299 ( .IN1(n2280), .IN2(keyinput30), .Q(n2279) );
  NAND2X0 U2300 ( .IN1(n2187), .IN2(n2281), .QN(n2280) );
  NAND3X0 U2301 ( .IN1(n2282), .IN2(n2283), .IN3(n2284), .QN(n2281) );
  AO21X1 U2302 ( .IN1(n2282), .IN2(n2283), .IN3(n2284), .Q(n2187) );
  NAND2X0 U2303 ( .IN1(n2196), .IN2(n2285), .QN(n2284) );
  NAND3X0 U2304 ( .IN1(N511), .IN2(n2286), .IN3(N18), .QN(n2285) );
  AO21X1 U2305 ( .IN1(N18), .IN2(N511), .IN3(n2286), .Q(n2196) );
  NAND2X0 U2306 ( .IN1(n2194), .IN2(n2287), .QN(n2286) );
  NAND3X0 U2307 ( .IN1(n2288), .IN2(n2289), .IN3(n2290), .QN(n2287) );
  AO21X1 U2308 ( .IN1(n2288), .IN2(n2289), .IN3(n2290), .Q(n2194) );
  NAND2X0 U2309 ( .IN1(n2202), .IN2(n2291), .QN(n2290) );
  NAND3X0 U2310 ( .IN1(N494), .IN2(n2292), .IN3(N35), .QN(n2291) );
  AO21X1 U2311 ( .IN1(N35), .IN2(N494), .IN3(n2292), .Q(n2202) );
  NAND2X0 U2312 ( .IN1(n2203), .IN2(n2293), .QN(n2292) );
  NAND3X0 U2313 ( .IN1(n2294), .IN2(n2295), .IN3(n2296), .QN(n2293) );
  AO21X1 U2314 ( .IN1(n2294), .IN2(n2295), .IN3(n2296), .Q(n2203) );
  NAND2X0 U2315 ( .IN1(n2208), .IN2(n2297), .QN(n2296) );
  NAND3X0 U2316 ( .IN1(N477), .IN2(n2298), .IN3(N52), .QN(n2297) );
  AO21X1 U2317 ( .IN1(N52), .IN2(N477), .IN3(n2298), .Q(n2208) );
  NAND2X0 U2318 ( .IN1(n2209), .IN2(n2299), .QN(n2298) );
  NAND3X0 U2319 ( .IN1(n2300), .IN2(n2301), .IN3(n2302), .QN(n2299) );
  AO21X1 U2320 ( .IN1(n2300), .IN2(n2301), .IN3(n2302), .Q(n2209) );
  AO21X1 U2321 ( .IN1(n2303), .IN2(n2304), .IN3(n2305), .Q(n2302) );
  INVX0 U2322 ( .INP(n2216), .ZN(n2305) );
  XNOR2X1 U2323 ( .IN1(n2306), .IN2(keyinput19), .Q(n2216) );
  OR2X1 U2324 ( .IN1(n2304), .IN2(n2303), .Q(n2306) );
  NAND2X0 U2325 ( .IN1(n2215), .IN2(n2307), .QN(n2304) );
  NAND3X0 U2326 ( .IN1(n2308), .IN2(n2309), .IN3(n2310), .QN(n2307) );
  AO21X1 U2327 ( .IN1(n2308), .IN2(n2309), .IN3(n2310), .Q(n2215) );
  NAND2X0 U2328 ( .IN1(n2220), .IN2(n2311), .QN(n2310) );
  NAND3X0 U2329 ( .IN1(N443), .IN2(n2312), .IN3(N86), .QN(n2311) );
  AO21X1 U2330 ( .IN1(N86), .IN2(N443), .IN3(n2312), .Q(n2220) );
  NAND2X0 U2331 ( .IN1(n2221), .IN2(n2313), .QN(n2312) );
  NAND3X0 U2332 ( .IN1(n2314), .IN2(n2315), .IN3(n2316), .QN(n2313) );
  AO21X1 U2333 ( .IN1(n2314), .IN2(n2315), .IN3(n2316), .Q(n2221) );
  NAND2X0 U2334 ( .IN1(n2226), .IN2(n2317), .QN(n2316) );
  NAND3X0 U2335 ( .IN1(N426), .IN2(n2318), .IN3(N103), .QN(n2317) );
  AO21X1 U2336 ( .IN1(N103), .IN2(N426), .IN3(n2318), .Q(n2226) );
  NAND2X0 U2337 ( .IN1(n2227), .IN2(n2319), .QN(n2318) );
  NAND3X0 U2338 ( .IN1(n2320), .IN2(n2321), .IN3(n2322), .QN(n2319) );
  AO21X1 U2339 ( .IN1(n2320), .IN2(n2321), .IN3(n2322), .Q(n2227) );
  NAND2X0 U2340 ( .IN1(n2232), .IN2(n2323), .QN(n2322) );
  NAND3X0 U2341 ( .IN1(N409), .IN2(n2324), .IN3(N120), .QN(n2323) );
  AO21X1 U2342 ( .IN1(N120), .IN2(N409), .IN3(n2324), .Q(n2232) );
  NAND2X0 U2343 ( .IN1(n2233), .IN2(n2325), .QN(n2324) );
  NAND3X0 U2344 ( .IN1(n2326), .IN2(n2327), .IN3(n2328), .QN(n2325) );
  AO21X1 U2345 ( .IN1(n2326), .IN2(n2327), .IN3(n2328), .Q(n2233) );
  NAND2X0 U2346 ( .IN1(n2238), .IN2(n2329), .QN(n2328) );
  NAND3X0 U2347 ( .IN1(N392), .IN2(n2330), .IN3(N137), .QN(n2329) );
  AO21X1 U2348 ( .IN1(N137), .IN2(N392), .IN3(n2330), .Q(n2238) );
  NAND2X0 U2349 ( .IN1(n2239), .IN2(n2331), .QN(n2330) );
  NAND3X0 U2350 ( .IN1(n2332), .IN2(n2333), .IN3(n2334), .QN(n2331) );
  AO21X1 U2351 ( .IN1(n2332), .IN2(n2333), .IN3(n2334), .Q(n2239) );
  NAND2X0 U2352 ( .IN1(n2244), .IN2(n2335), .QN(n2334) );
  NAND3X0 U2353 ( .IN1(N375), .IN2(n2336), .IN3(N154), .QN(n2335) );
  AO21X1 U2354 ( .IN1(N154), .IN2(N375), .IN3(n2336), .Q(n2244) );
  NAND2X0 U2355 ( .IN1(n2245), .IN2(n2337), .QN(n2336) );
  NAND3X0 U2356 ( .IN1(n2338), .IN2(n2339), .IN3(n2340), .QN(n2337) );
  AO21X1 U2357 ( .IN1(n2338), .IN2(n2339), .IN3(n2340), .Q(n2245) );
  NAND2X0 U2358 ( .IN1(n2250), .IN2(n2341), .QN(n2340) );
  NAND3X0 U2359 ( .IN1(N358), .IN2(n2342), .IN3(N171), .QN(n2341) );
  AO21X1 U2360 ( .IN1(N171), .IN2(N358), .IN3(n2342), .Q(n2250) );
  NAND2X0 U2361 ( .IN1(n2251), .IN2(n2343), .QN(n2342) );
  NAND3X0 U2362 ( .IN1(n2344), .IN2(n2345), .IN3(n2346), .QN(n2343) );
  AO21X1 U2363 ( .IN1(n2344), .IN2(n2345), .IN3(n2346), .Q(n2251) );
  NAND2X0 U2364 ( .IN1(n2256), .IN2(n2347), .QN(n2346) );
  NAND3X0 U2365 ( .IN1(N341), .IN2(n2348), .IN3(N188), .QN(n2347) );
  AO21X1 U2366 ( .IN1(N188), .IN2(N341), .IN3(n2348), .Q(n2256) );
  NAND2X0 U2367 ( .IN1(n2257), .IN2(n2349), .QN(n2348) );
  NAND3X0 U2368 ( .IN1(n2350), .IN2(n2351), .IN3(n2352), .QN(n2349) );
  AO21X1 U2369 ( .IN1(n2350), .IN2(n2351), .IN3(n2352), .Q(n2257) );
  NAND2X0 U2370 ( .IN1(n2262), .IN2(n2353), .QN(n2352) );
  NAND3X0 U2371 ( .IN1(N324), .IN2(n2354), .IN3(N205), .QN(n2353) );
  AO21X1 U2372 ( .IN1(N205), .IN2(N324), .IN3(n2354), .Q(n2262) );
  NAND2X0 U2373 ( .IN1(n2263), .IN2(n2355), .QN(n2354) );
  NAND3X0 U2374 ( .IN1(n2356), .IN2(n2357), .IN3(n2358), .QN(n2355) );
  AO21X1 U2375 ( .IN1(n2356), .IN2(n2357), .IN3(n2358), .Q(n2263) );
  NAND2X0 U2376 ( .IN1(n2271), .IN2(n2359), .QN(n2358) );
  NAND3X0 U2377 ( .IN1(N307), .IN2(n2360), .IN3(N222), .QN(n2359) );
  AO21X1 U2378 ( .IN1(N222), .IN2(N307), .IN3(n2360), .Q(n2271) );
  NAND2X0 U2379 ( .IN1(n2272), .IN2(n2361), .QN(n2360) );
  NAND3X0 U2380 ( .IN1(n2362), .IN2(n2274), .IN3(n2363), .QN(n2361) );
  AO21X1 U2381 ( .IN1(n2362), .IN2(n2274), .IN3(n2363), .Q(n2272) );
  NAND3X0 U2382 ( .IN1(N256), .IN2(N239), .IN3(n2364), .QN(n2274) );
  AO22X1 U2383 ( .IN1(N290), .IN2(N239), .IN3(N273), .IN4(N256), .Q(n2362) );
  AND2X1 U2384 ( .IN1(N69), .IN2(N460), .Q(n2303) );
  NAND2X0 U2385 ( .IN1(n2282), .IN2(n2365), .QN(N5971) );
  NAND3X0 U2386 ( .IN1(N511), .IN2(n2366), .IN3(N1), .QN(n2365) );
  AO21X1 U2387 ( .IN1(N1), .IN2(N511), .IN3(n2366), .Q(n2282) );
  NAND2X0 U2388 ( .IN1(n2283), .IN2(n2367), .QN(n2366) );
  NAND3X0 U2389 ( .IN1(n2368), .IN2(n2369), .IN3(n2370), .QN(n2367) );
  AO21X1 U2390 ( .IN1(n2368), .IN2(n2369), .IN3(n2370), .Q(n2283) );
  NAND2X0 U2391 ( .IN1(n2288), .IN2(n2371), .QN(n2370) );
  NAND3X0 U2392 ( .IN1(N494), .IN2(n2372), .IN3(N18), .QN(n2371) );
  AO21X1 U2393 ( .IN1(N18), .IN2(N494), .IN3(n2372), .Q(n2288) );
  NAND2X0 U2394 ( .IN1(n2289), .IN2(n2373), .QN(n2372) );
  NAND3X0 U2395 ( .IN1(n2374), .IN2(n2375), .IN3(n2376), .QN(n2373) );
  AO21X1 U2396 ( .IN1(n2374), .IN2(n2375), .IN3(n2376), .Q(n2289) );
  NAND2X0 U2397 ( .IN1(n2294), .IN2(n2377), .QN(n2376) );
  NAND3X0 U2398 ( .IN1(N477), .IN2(n2378), .IN3(N35), .QN(n2377) );
  AO21X1 U2399 ( .IN1(N35), .IN2(N477), .IN3(n2378), .Q(n2294) );
  NAND2X0 U2400 ( .IN1(n2295), .IN2(n2379), .QN(n2378) );
  NAND3X0 U2401 ( .IN1(n2380), .IN2(n2381), .IN3(n2382), .QN(n2379) );
  AO21X1 U2402 ( .IN1(n2380), .IN2(n2381), .IN3(n2382), .Q(n2295) );
  NAND2X0 U2403 ( .IN1(n2300), .IN2(n2383), .QN(n2382) );
  NAND3X0 U2404 ( .IN1(N460), .IN2(n2384), .IN3(N52), .QN(n2383) );
  AO21X1 U2405 ( .IN1(N52), .IN2(N460), .IN3(n2384), .Q(n2300) );
  NAND2X0 U2406 ( .IN1(n2301), .IN2(n2385), .QN(n2384) );
  NAND3X0 U2407 ( .IN1(n2386), .IN2(n2387), .IN3(n2388), .QN(n2385) );
  AO21X1 U2408 ( .IN1(n2386), .IN2(n2387), .IN3(n2388), .Q(n2301) );
  NAND2X0 U2409 ( .IN1(n2308), .IN2(n2389), .QN(n2388) );
  NAND3X0 U2410 ( .IN1(N443), .IN2(n2390), .IN3(N69), .QN(n2389) );
  AO21X1 U2411 ( .IN1(N69), .IN2(N443), .IN3(n2390), .Q(n2308) );
  NAND2X0 U2412 ( .IN1(n2309), .IN2(n2391), .QN(n2390) );
  NAND3X0 U2413 ( .IN1(n2392), .IN2(n2393), .IN3(n2394), .QN(n2391) );
  AO21X1 U2414 ( .IN1(n2392), .IN2(n2393), .IN3(n2394), .Q(n2309) );
  XNOR2X1 U2415 ( .IN1(n2395), .IN2(keyinput16), .Q(n2394) );
  NAND2X0 U2416 ( .IN1(n2314), .IN2(n2396), .QN(n2395) );
  NAND3X0 U2417 ( .IN1(N426), .IN2(n2397), .IN3(N86), .QN(n2396) );
  AO21X1 U2418 ( .IN1(N86), .IN2(N426), .IN3(n2397), .Q(n2314) );
  NAND2X0 U2419 ( .IN1(n2315), .IN2(n2398), .QN(n2397) );
  NAND3X0 U2420 ( .IN1(n2399), .IN2(n2400), .IN3(n2401), .QN(n2398) );
  AO21X1 U2421 ( .IN1(n2399), .IN2(n2400), .IN3(n2401), .Q(n2315) );
  NAND2X0 U2422 ( .IN1(n2320), .IN2(n2402), .QN(n2401) );
  NAND3X0 U2423 ( .IN1(N409), .IN2(n2403), .IN3(N103), .QN(n2402) );
  AO21X1 U2424 ( .IN1(N103), .IN2(N409), .IN3(n2403), .Q(n2320) );
  NAND2X0 U2425 ( .IN1(n2321), .IN2(n2404), .QN(n2403) );
  NAND3X0 U2426 ( .IN1(n2405), .IN2(n2406), .IN3(n2407), .QN(n2404) );
  AO21X1 U2427 ( .IN1(n2405), .IN2(n2406), .IN3(n2407), .Q(n2321) );
  NAND2X0 U2428 ( .IN1(n2326), .IN2(n2408), .QN(n2407) );
  NAND3X0 U2429 ( .IN1(N392), .IN2(n2409), .IN3(N120), .QN(n2408) );
  AO21X1 U2430 ( .IN1(N120), .IN2(N392), .IN3(n2409), .Q(n2326) );
  NAND2X0 U2431 ( .IN1(n2327), .IN2(n2410), .QN(n2409) );
  NAND3X0 U2432 ( .IN1(n2411), .IN2(n2412), .IN3(n2413), .QN(n2410) );
  AO21X1 U2433 ( .IN1(n2411), .IN2(n2412), .IN3(n2413), .Q(n2327) );
  NAND2X0 U2434 ( .IN1(n2332), .IN2(n2414), .QN(n2413) );
  NAND3X0 U2435 ( .IN1(N375), .IN2(n2415), .IN3(N137), .QN(n2414) );
  AO21X1 U2436 ( .IN1(N137), .IN2(N375), .IN3(n2415), .Q(n2332) );
  NAND2X0 U2437 ( .IN1(n2333), .IN2(n2416), .QN(n2415) );
  NAND3X0 U2438 ( .IN1(n2417), .IN2(n2418), .IN3(n2419), .QN(n2416) );
  AO21X1 U2439 ( .IN1(n2417), .IN2(n2418), .IN3(n2419), .Q(n2333) );
  NAND2X0 U2440 ( .IN1(n2338), .IN2(n2420), .QN(n2419) );
  NAND3X0 U2441 ( .IN1(N358), .IN2(n2421), .IN3(N154), .QN(n2420) );
  AO21X1 U2442 ( .IN1(N154), .IN2(N358), .IN3(n2421), .Q(n2338) );
  NAND2X0 U2443 ( .IN1(n2339), .IN2(n2422), .QN(n2421) );
  NAND3X0 U2444 ( .IN1(n2423), .IN2(n2424), .IN3(n2425), .QN(n2422) );
  AO21X1 U2445 ( .IN1(n2423), .IN2(n2424), .IN3(n2425), .Q(n2339) );
  NAND2X0 U2446 ( .IN1(n2344), .IN2(n2426), .QN(n2425) );
  NAND3X0 U2447 ( .IN1(N341), .IN2(n2427), .IN3(N171), .QN(n2426) );
  AO21X1 U2448 ( .IN1(N171), .IN2(N341), .IN3(n2427), .Q(n2344) );
  NAND2X0 U2449 ( .IN1(n2345), .IN2(n2428), .QN(n2427) );
  NAND3X0 U2450 ( .IN1(n2429), .IN2(n2430), .IN3(n2431), .QN(n2428) );
  AO21X1 U2451 ( .IN1(n2429), .IN2(n2430), .IN3(n2431), .Q(n2345) );
  NAND2X0 U2452 ( .IN1(n2350), .IN2(n2432), .QN(n2431) );
  NAND3X0 U2453 ( .IN1(N324), .IN2(n2433), .IN3(N188), .QN(n2432) );
  AO21X1 U2454 ( .IN1(N188), .IN2(N324), .IN3(n2433), .Q(n2350) );
  NAND2X0 U2455 ( .IN1(n2351), .IN2(n2434), .QN(n2433) );
  NAND3X0 U2456 ( .IN1(n2435), .IN2(n2436), .IN3(n2437), .QN(n2434) );
  AO21X1 U2457 ( .IN1(n2435), .IN2(n2436), .IN3(n2437), .Q(n2351) );
  NAND2X0 U2458 ( .IN1(n2356), .IN2(n2438), .QN(n2437) );
  NAND4X0 U2459 ( .IN1(N205), .IN2(N307), .IN3(n2439), .IN4(n2440), .QN(n2438)
         );
  AO22X1 U2460 ( .IN1(N205), .IN2(N307), .IN3(n2439), .IN4(n2440), .Q(n2356)
         );
  NAND2X0 U2461 ( .IN1(n2363), .IN2(n2357), .QN(n2440) );
  XNOR2X1 U2462 ( .IN1(n2441), .IN2(keyinput5), .Q(n2439) );
  NAND2X0 U2463 ( .IN1(n2442), .IN2(n2357), .QN(n2441) );
  AO21X1 U2464 ( .IN1(n2443), .IN2(n2444), .IN3(n2445), .Q(n2357) );
  INVX0 U2465 ( .INP(n2363), .ZN(n2444) );
  NOR2X0 U2466 ( .IN1(n2446), .IN2(n2447), .QN(n2363) );
  AO21X1 U2467 ( .IN1(N222), .IN2(N290), .IN3(n2447), .Q(n2443) );
  MUX21X1 U2468 ( .IN1(n2448), .IN2(n2449), .S(keyinput3), .Q(n2447) );
  AOI21X1 U2469 ( .IN1(N290), .IN2(N222), .IN3(n2446), .QN(n2449) );
  NAND2X0 U2470 ( .IN1(N273), .IN2(N239), .QN(n2446) );
  NAND2X0 U2471 ( .IN1(N239), .IN2(n2450), .QN(n2448) );
  OAI21X1 U2472 ( .IN1(n2451), .IN2(N222), .IN3(n2452), .QN(n2450) );
  INVX0 U2473 ( .INP(n2453), .ZN(n2412) );
  NAND2X0 U2474 ( .IN1(n2368), .IN2(n2454), .QN(N5672) );
  NAND3X0 U2475 ( .IN1(N494), .IN2(n2455), .IN3(N1), .QN(n2454) );
  AO21X1 U2476 ( .IN1(N1), .IN2(N494), .IN3(n2455), .Q(n2368) );
  NAND2X0 U2477 ( .IN1(n2369), .IN2(n2456), .QN(n2455) );
  NAND3X0 U2478 ( .IN1(n2457), .IN2(n2458), .IN3(n2459), .QN(n2456) );
  AO21X1 U2479 ( .IN1(n2457), .IN2(n2458), .IN3(n2459), .Q(n2369) );
  NAND2X0 U2480 ( .IN1(n2374), .IN2(n2460), .QN(n2459) );
  NAND3X0 U2481 ( .IN1(N477), .IN2(n2461), .IN3(N18), .QN(n2460) );
  AO21X1 U2482 ( .IN1(N18), .IN2(N477), .IN3(n2461), .Q(n2374) );
  NAND2X0 U2483 ( .IN1(n2375), .IN2(n2462), .QN(n2461) );
  NAND3X0 U2484 ( .IN1(n2463), .IN2(n2464), .IN3(n2465), .QN(n2462) );
  AO21X1 U2485 ( .IN1(n2463), .IN2(n2464), .IN3(n2465), .Q(n2375) );
  NAND2X0 U2486 ( .IN1(n2380), .IN2(n2466), .QN(n2465) );
  NAND3X0 U2487 ( .IN1(N460), .IN2(n2467), .IN3(N35), .QN(n2466) );
  AO21X1 U2488 ( .IN1(N35), .IN2(N460), .IN3(n2467), .Q(n2380) );
  NAND2X0 U2489 ( .IN1(n2381), .IN2(n2468), .QN(n2467) );
  NAND3X0 U2490 ( .IN1(n2469), .IN2(n2470), .IN3(n2471), .QN(n2468) );
  AO21X1 U2491 ( .IN1(n2469), .IN2(n2470), .IN3(n2471), .Q(n2381) );
  NAND2X0 U2492 ( .IN1(n2386), .IN2(n2472), .QN(n2471) );
  NAND3X0 U2493 ( .IN1(N443), .IN2(n2473), .IN3(N52), .QN(n2472) );
  AO21X1 U2494 ( .IN1(N52), .IN2(N443), .IN3(n2473), .Q(n2386) );
  NAND2X0 U2495 ( .IN1(n2387), .IN2(n2474), .QN(n2473) );
  NAND3X0 U2496 ( .IN1(n2475), .IN2(n2476), .IN3(n2477), .QN(n2474) );
  AO21X1 U2497 ( .IN1(n2477), .IN2(n2476), .IN3(n2475), .Q(n2387) );
  NAND2X0 U2498 ( .IN1(n2392), .IN2(n2478), .QN(n2475) );
  NAND3X0 U2499 ( .IN1(N426), .IN2(n2479), .IN3(N69), .QN(n2478) );
  AO21X1 U2500 ( .IN1(N69), .IN2(N426), .IN3(n2479), .Q(n2392) );
  NAND2X0 U2501 ( .IN1(n2393), .IN2(n2480), .QN(n2479) );
  NAND3X0 U2502 ( .IN1(n2481), .IN2(n2482), .IN3(n2483), .QN(n2480) );
  AO21X1 U2503 ( .IN1(n2481), .IN2(n2482), .IN3(n2483), .Q(n2393) );
  NAND2X0 U2504 ( .IN1(n2399), .IN2(n2484), .QN(n2483) );
  NAND3X0 U2505 ( .IN1(N409), .IN2(n2485), .IN3(N86), .QN(n2484) );
  AO21X1 U2506 ( .IN1(N86), .IN2(N409), .IN3(n2485), .Q(n2399) );
  NAND2X0 U2507 ( .IN1(n2400), .IN2(n2486), .QN(n2485) );
  NAND3X0 U2508 ( .IN1(n2487), .IN2(n2488), .IN3(n2489), .QN(n2486) );
  AO21X1 U2509 ( .IN1(n2487), .IN2(n2488), .IN3(n2489), .Q(n2400) );
  NAND2X0 U2510 ( .IN1(n2405), .IN2(n2490), .QN(n2489) );
  NAND3X0 U2511 ( .IN1(N392), .IN2(n2491), .IN3(N103), .QN(n2490) );
  AO21X1 U2512 ( .IN1(N103), .IN2(N392), .IN3(n2491), .Q(n2405) );
  NAND2X0 U2513 ( .IN1(n2406), .IN2(n2492), .QN(n2491) );
  NAND3X0 U2514 ( .IN1(n2493), .IN2(n2494), .IN3(n2495), .QN(n2492) );
  AO21X1 U2515 ( .IN1(n2493), .IN2(n2494), .IN3(n2495), .Q(n2406) );
  NAND2X0 U2516 ( .IN1(n2411), .IN2(n2496), .QN(n2495) );
  NAND3X0 U2517 ( .IN1(N375), .IN2(n2497), .IN3(N120), .QN(n2496) );
  AO21X1 U2518 ( .IN1(N120), .IN2(N375), .IN3(n2497), .Q(n2411) );
  AO21X1 U2519 ( .IN1(n2498), .IN2(n2499), .IN3(n2453), .Q(n2497) );
  NOR2X0 U2520 ( .IN1(n2499), .IN2(n2498), .QN(n2453) );
  NAND2X0 U2521 ( .IN1(n2417), .IN2(n2500), .QN(n2499) );
  NAND3X0 U2522 ( .IN1(N358), .IN2(n2501), .IN3(N137), .QN(n2500) );
  AO21X1 U2523 ( .IN1(N137), .IN2(N358), .IN3(n2501), .Q(n2417) );
  NAND2X0 U2524 ( .IN1(n2418), .IN2(n2502), .QN(n2501) );
  NAND3X0 U2525 ( .IN1(n2503), .IN2(n2504), .IN3(n2505), .QN(n2502) );
  AO21X1 U2526 ( .IN1(n2503), .IN2(n2504), .IN3(n2505), .Q(n2418) );
  NAND2X0 U2527 ( .IN1(n2423), .IN2(n2506), .QN(n2505) );
  NAND3X0 U2528 ( .IN1(N341), .IN2(n2507), .IN3(N154), .QN(n2506) );
  AO21X1 U2529 ( .IN1(N154), .IN2(N341), .IN3(n2507), .Q(n2423) );
  NAND2X0 U2530 ( .IN1(n2424), .IN2(n2508), .QN(n2507) );
  NAND3X0 U2531 ( .IN1(n2509), .IN2(n2510), .IN3(n2511), .QN(n2508) );
  AO21X1 U2532 ( .IN1(n2509), .IN2(n2510), .IN3(n2511), .Q(n2424) );
  NAND2X0 U2533 ( .IN1(n2429), .IN2(n2512), .QN(n2511) );
  NAND3X0 U2534 ( .IN1(N324), .IN2(n2513), .IN3(N171), .QN(n2512) );
  AO21X1 U2535 ( .IN1(N171), .IN2(N324), .IN3(n2513), .Q(n2429) );
  NAND2X0 U2536 ( .IN1(n2430), .IN2(n2514), .QN(n2513) );
  NAND3X0 U2537 ( .IN1(n2515), .IN2(n2516), .IN3(n2517), .QN(n2514) );
  AO21X1 U2538 ( .IN1(n2515), .IN2(n2516), .IN3(n2517), .Q(n2430) );
  NAND2X0 U2539 ( .IN1(n2435), .IN2(n2518), .QN(n2517) );
  NAND3X0 U2540 ( .IN1(N307), .IN2(n2519), .IN3(N188), .QN(n2518) );
  AO21X1 U2541 ( .IN1(N188), .IN2(N307), .IN3(n2519), .Q(n2435) );
  OAI21X1 U2542 ( .IN1(n2520), .IN2(n2445), .IN3(n2436), .QN(n2519) );
  AO21X1 U2543 ( .IN1(n2521), .IN2(n2442), .IN3(n2522), .Q(n2436) );
  AO22X1 U2544 ( .IN1(N205), .IN2(N290), .IN3(N222), .IN4(N273), .Q(n2521) );
  INVX0 U2545 ( .INP(n2442), .ZN(n2445) );
  NAND3X0 U2546 ( .IN1(N222), .IN2(n2364), .IN3(N205), .QN(n2442) );
  INVX0 U2547 ( .INP(n2523), .ZN(n2477) );
  NAND2X0 U2548 ( .IN1(n2457), .IN2(n2524), .QN(N5308) );
  NAND3X0 U2549 ( .IN1(N477), .IN2(n2525), .IN3(N1), .QN(n2524) );
  AO21X1 U2550 ( .IN1(N1), .IN2(N477), .IN3(n2525), .Q(n2457) );
  NAND2X0 U2551 ( .IN1(n2458), .IN2(n2526), .QN(n2525) );
  NAND3X0 U2552 ( .IN1(n2527), .IN2(n2528), .IN3(n2529), .QN(n2526) );
  AO21X1 U2553 ( .IN1(n2527), .IN2(n2528), .IN3(n2529), .Q(n2458) );
  NAND2X0 U2554 ( .IN1(n2463), .IN2(n2530), .QN(n2529) );
  NAND3X0 U2555 ( .IN1(N460), .IN2(n2531), .IN3(N18), .QN(n2530) );
  AO21X1 U2556 ( .IN1(N18), .IN2(N460), .IN3(n2531), .Q(n2463) );
  NAND2X0 U2557 ( .IN1(n2464), .IN2(n2532), .QN(n2531) );
  NAND3X0 U2558 ( .IN1(n2533), .IN2(n2534), .IN3(n2535), .QN(n2532) );
  AO21X1 U2559 ( .IN1(n2533), .IN2(n2534), .IN3(n2535), .Q(n2464) );
  NAND2X0 U2560 ( .IN1(n2469), .IN2(n2536), .QN(n2535) );
  NAND3X0 U2561 ( .IN1(N443), .IN2(n2537), .IN3(N35), .QN(n2536) );
  AO21X1 U2562 ( .IN1(N35), .IN2(N443), .IN3(n2537), .Q(n2469) );
  NAND2X0 U2563 ( .IN1(n2470), .IN2(n2538), .QN(n2537) );
  NAND3X0 U2564 ( .IN1(n2539), .IN2(n2540), .IN3(n2541), .QN(n2538) );
  AO21X1 U2565 ( .IN1(n2539), .IN2(n2540), .IN3(n2541), .Q(n2470) );
  AO21X1 U2566 ( .IN1(n2542), .IN2(n2543), .IN3(n2523), .Q(n2541) );
  NOR2X0 U2567 ( .IN1(n2543), .IN2(n2542), .QN(n2523) );
  NAND2X0 U2568 ( .IN1(n2476), .IN2(n2544), .QN(n2543) );
  NAND3X0 U2569 ( .IN1(n2545), .IN2(n2546), .IN3(n2547), .QN(n2544) );
  AO21X1 U2570 ( .IN1(n2545), .IN2(n2546), .IN3(n2547), .Q(n2476) );
  NAND2X0 U2571 ( .IN1(n2481), .IN2(n2548), .QN(n2547) );
  NAND3X0 U2572 ( .IN1(N409), .IN2(n2549), .IN3(N69), .QN(n2548) );
  AO21X1 U2573 ( .IN1(N69), .IN2(N409), .IN3(n2549), .Q(n2481) );
  NAND2X0 U2574 ( .IN1(n2482), .IN2(n2550), .QN(n2549) );
  NAND3X0 U2575 ( .IN1(n2551), .IN2(n2552), .IN3(n2553), .QN(n2550) );
  AO21X1 U2576 ( .IN1(n2551), .IN2(n2552), .IN3(n2553), .Q(n2482) );
  NAND2X0 U2577 ( .IN1(n2487), .IN2(n2554), .QN(n2553) );
  NAND3X0 U2578 ( .IN1(N392), .IN2(n2555), .IN3(N86), .QN(n2554) );
  AO21X1 U2579 ( .IN1(N86), .IN2(N392), .IN3(n2555), .Q(n2487) );
  NAND2X0 U2580 ( .IN1(n2488), .IN2(n2556), .QN(n2555) );
  NAND3X0 U2581 ( .IN1(n2557), .IN2(n2558), .IN3(n2559), .QN(n2556) );
  AO21X1 U2582 ( .IN1(n2557), .IN2(n2558), .IN3(n2559), .Q(n2488) );
  NAND2X0 U2583 ( .IN1(n2493), .IN2(n2560), .QN(n2559) );
  NAND3X0 U2584 ( .IN1(N375), .IN2(n2561), .IN3(N103), .QN(n2560) );
  AO21X1 U2585 ( .IN1(N103), .IN2(N375), .IN3(n2561), .Q(n2493) );
  NAND2X0 U2586 ( .IN1(n2494), .IN2(n2562), .QN(n2561) );
  NAND4X0 U2587 ( .IN1(n2563), .IN2(n2564), .IN3(n2565), .IN4(n2566), .QN(
        n2562) );
  AO22X1 U2588 ( .IN1(n2565), .IN2(n2566), .IN3(n2563), .IN4(n2564), .Q(n2494)
         );
  AO21X1 U2589 ( .IN1(N120), .IN2(N358), .IN3(n2567), .Q(n2564) );
  INVX0 U2590 ( .INP(n2568), .ZN(n2567) );
  XOR2X1 U2591 ( .IN1(n2569), .IN2(keyinput12), .Q(n2563) );
  NAND2X0 U2592 ( .IN1(n2498), .IN2(n2570), .QN(n2569) );
  AND2X1 U2593 ( .IN1(n2568), .IN2(n2571), .Q(n2498) );
  NAND3X0 U2594 ( .IN1(n2570), .IN2(n2571), .IN3(n2572), .QN(n2568) );
  NAND2X0 U2595 ( .IN1(N120), .IN2(N358), .QN(n2572) );
  AO21X1 U2596 ( .IN1(n2573), .IN2(n2574), .IN3(n2575), .Q(n2571) );
  NAND3X0 U2597 ( .IN1(n2573), .IN2(n2574), .IN3(n2575), .QN(n2570) );
  NAND2X0 U2598 ( .IN1(n2503), .IN2(n2576), .QN(n2575) );
  NAND3X0 U2599 ( .IN1(N341), .IN2(n2577), .IN3(N137), .QN(n2576) );
  AO21X1 U2600 ( .IN1(N137), .IN2(N341), .IN3(n2577), .Q(n2503) );
  NAND2X0 U2601 ( .IN1(n2504), .IN2(n2578), .QN(n2577) );
  NAND3X0 U2602 ( .IN1(n2579), .IN2(n2580), .IN3(n2581), .QN(n2578) );
  AO21X1 U2603 ( .IN1(n2579), .IN2(n2580), .IN3(n2581), .Q(n2504) );
  NAND2X0 U2604 ( .IN1(n2509), .IN2(n2582), .QN(n2581) );
  NAND3X0 U2605 ( .IN1(N324), .IN2(n2583), .IN3(N154), .QN(n2582) );
  AO21X1 U2606 ( .IN1(N154), .IN2(N324), .IN3(n2583), .Q(n2509) );
  NAND2X0 U2607 ( .IN1(n2510), .IN2(n2584), .QN(n2583) );
  NAND3X0 U2608 ( .IN1(n2585), .IN2(n2586), .IN3(n2587), .QN(n2584) );
  AO21X1 U2609 ( .IN1(n2585), .IN2(n2586), .IN3(n2587), .Q(n2510) );
  NAND2X0 U2610 ( .IN1(n2515), .IN2(n2588), .QN(n2587) );
  NAND3X0 U2611 ( .IN1(N307), .IN2(n2589), .IN3(N171), .QN(n2588) );
  AO21X1 U2612 ( .IN1(N171), .IN2(N307), .IN3(n2589), .Q(n2515) );
  OAI21X1 U2613 ( .IN1(n2590), .IN2(n2522), .IN3(n2516), .QN(n2589) );
  AO21X1 U2614 ( .IN1(n2591), .IN2(n2520), .IN3(n2592), .Q(n2516) );
  AO22X1 U2615 ( .IN1(N188), .IN2(N290), .IN3(N205), .IN4(N273), .Q(n2591) );
  INVX0 U2616 ( .INP(n2520), .ZN(n2522) );
  NAND3X0 U2617 ( .IN1(N205), .IN2(n2364), .IN3(N188), .QN(n2520) );
  XOR2X1 U2618 ( .IN1(n2593), .IN2(keyinput0), .Q(n2542) );
  NAND2X0 U2619 ( .IN1(N52), .IN2(N426), .QN(n2593) );
  NAND2X0 U2620 ( .IN1(n2527), .IN2(n2594), .QN(N4946) );
  NAND3X0 U2621 ( .IN1(N460), .IN2(n2595), .IN3(N1), .QN(n2594) );
  AO21X1 U2622 ( .IN1(N1), .IN2(N460), .IN3(n2595), .Q(n2527) );
  NAND2X0 U2623 ( .IN1(n2528), .IN2(n2596), .QN(n2595) );
  NAND3X0 U2624 ( .IN1(n2597), .IN2(n2598), .IN3(n2599), .QN(n2596) );
  AO21X1 U2625 ( .IN1(n2597), .IN2(n2598), .IN3(n2599), .Q(n2528) );
  NAND2X0 U2626 ( .IN1(n2533), .IN2(n2600), .QN(n2599) );
  NAND3X0 U2627 ( .IN1(N443), .IN2(n2601), .IN3(N18), .QN(n2600) );
  AO21X1 U2628 ( .IN1(N18), .IN2(N443), .IN3(n2601), .Q(n2533) );
  NAND2X0 U2629 ( .IN1(n2534), .IN2(n2602), .QN(n2601) );
  NAND3X0 U2630 ( .IN1(n2603), .IN2(n2604), .IN3(n2605), .QN(n2602) );
  AO21X1 U2631 ( .IN1(n2603), .IN2(n2604), .IN3(n2605), .Q(n2534) );
  NAND2X0 U2632 ( .IN1(n2539), .IN2(n2606), .QN(n2605) );
  NAND3X0 U2633 ( .IN1(N426), .IN2(n2607), .IN3(N35), .QN(n2606) );
  AO21X1 U2634 ( .IN1(N35), .IN2(N426), .IN3(n2607), .Q(n2539) );
  NAND2X0 U2635 ( .IN1(n2540), .IN2(n2608), .QN(n2607) );
  NAND3X0 U2636 ( .IN1(n2609), .IN2(n2610), .IN3(n2611), .QN(n2608) );
  AO21X1 U2637 ( .IN1(n2609), .IN2(n2610), .IN3(n2611), .Q(n2540) );
  NAND2X0 U2638 ( .IN1(n2545), .IN2(n2612), .QN(n2611) );
  NAND3X0 U2639 ( .IN1(N409), .IN2(n2613), .IN3(N52), .QN(n2612) );
  AO21X1 U2640 ( .IN1(N52), .IN2(N409), .IN3(n2613), .Q(n2545) );
  NAND2X0 U2641 ( .IN1(n2546), .IN2(n2614), .QN(n2613) );
  NAND3X0 U2642 ( .IN1(n2615), .IN2(n2616), .IN3(n2617), .QN(n2614) );
  AO21X1 U2643 ( .IN1(n2615), .IN2(n2616), .IN3(n2617), .Q(n2546) );
  NAND2X0 U2644 ( .IN1(n2551), .IN2(n2618), .QN(n2617) );
  NAND3X0 U2645 ( .IN1(N392), .IN2(n2619), .IN3(N69), .QN(n2618) );
  AO21X1 U2646 ( .IN1(N69), .IN2(N392), .IN3(n2619), .Q(n2551) );
  NAND2X0 U2647 ( .IN1(n2552), .IN2(n2620), .QN(n2619) );
  NAND3X0 U2648 ( .IN1(n2621), .IN2(n2622), .IN3(n2623), .QN(n2620) );
  AO21X1 U2649 ( .IN1(n2621), .IN2(n2622), .IN3(n2623), .Q(n2552) );
  NAND2X0 U2650 ( .IN1(n2557), .IN2(n2624), .QN(n2623) );
  NAND3X0 U2651 ( .IN1(N375), .IN2(n2625), .IN3(N86), .QN(n2624) );
  AO21X1 U2652 ( .IN1(N86), .IN2(N375), .IN3(n2625), .Q(n2557) );
  NAND2X0 U2653 ( .IN1(n2558), .IN2(n2626), .QN(n2625) );
  NAND3X0 U2654 ( .IN1(n2627), .IN2(n2628), .IN3(n2629), .QN(n2626) );
  AO21X1 U2655 ( .IN1(n2627), .IN2(n2628), .IN3(n2629), .Q(n2558) );
  NAND2X0 U2656 ( .IN1(n2565), .IN2(n2630), .QN(n2629) );
  NAND3X0 U2657 ( .IN1(N358), .IN2(n2631), .IN3(N103), .QN(n2630) );
  AO21X1 U2658 ( .IN1(N103), .IN2(N358), .IN3(n2631), .Q(n2565) );
  NAND2X0 U2659 ( .IN1(n2566), .IN2(n2632), .QN(n2631) );
  NAND3X0 U2660 ( .IN1(n2633), .IN2(n2634), .IN3(n2635), .QN(n2632) );
  AO21X1 U2661 ( .IN1(n2633), .IN2(n2634), .IN3(n2635), .Q(n2566) );
  NAND2X0 U2662 ( .IN1(n2573), .IN2(n2636), .QN(n2635) );
  NAND3X0 U2663 ( .IN1(N341), .IN2(n2637), .IN3(N120), .QN(n2636) );
  AO21X1 U2664 ( .IN1(N120), .IN2(N341), .IN3(n2637), .Q(n2573) );
  NAND2X0 U2665 ( .IN1(n2574), .IN2(n2638), .QN(n2637) );
  NAND3X0 U2666 ( .IN1(n2639), .IN2(n2640), .IN3(n2641), .QN(n2638) );
  AO21X1 U2667 ( .IN1(n2639), .IN2(n2640), .IN3(n2641), .Q(n2574) );
  NAND2X0 U2668 ( .IN1(n2579), .IN2(n2642), .QN(n2641) );
  NAND3X0 U2669 ( .IN1(N324), .IN2(n2643), .IN3(N137), .QN(n2642) );
  AO21X1 U2670 ( .IN1(N137), .IN2(N324), .IN3(n2643), .Q(n2579) );
  NAND2X0 U2671 ( .IN1(n2580), .IN2(n2644), .QN(n2643) );
  NAND3X0 U2672 ( .IN1(n2645), .IN2(n2646), .IN3(n2647), .QN(n2644) );
  AO21X1 U2673 ( .IN1(n2645), .IN2(n2646), .IN3(n2647), .Q(n2580) );
  NAND2X0 U2674 ( .IN1(n2585), .IN2(n2648), .QN(n2647) );
  NAND3X0 U2675 ( .IN1(N307), .IN2(n2649), .IN3(N154), .QN(n2648) );
  AO21X1 U2676 ( .IN1(N154), .IN2(N307), .IN3(n2649), .Q(n2585) );
  OAI21X1 U2677 ( .IN1(n2650), .IN2(n2592), .IN3(n2586), .QN(n2649) );
  AO21X1 U2678 ( .IN1(n2651), .IN2(n2590), .IN3(n2652), .Q(n2586) );
  AO22X1 U2679 ( .IN1(N171), .IN2(N290), .IN3(N188), .IN4(N273), .Q(n2651) );
  INVX0 U2680 ( .INP(n2590), .ZN(n2592) );
  NAND3X0 U2681 ( .IN1(N188), .IN2(n2364), .IN3(N171), .QN(n2590) );
  NAND2X0 U2682 ( .IN1(n2597), .IN2(n2653), .QN(N4591) );
  NAND3X0 U2683 ( .IN1(N443), .IN2(n2654), .IN3(N1), .QN(n2653) );
  AO21X1 U2684 ( .IN1(N1), .IN2(N443), .IN3(n2654), .Q(n2597) );
  NAND2X0 U2685 ( .IN1(n2598), .IN2(n2655), .QN(n2654) );
  NAND3X0 U2686 ( .IN1(n2656), .IN2(n2657), .IN3(n2658), .QN(n2655) );
  AO21X1 U2687 ( .IN1(n2656), .IN2(n2657), .IN3(n2658), .Q(n2598) );
  NAND2X0 U2688 ( .IN1(n2603), .IN2(n2659), .QN(n2658) );
  NAND3X0 U2689 ( .IN1(N426), .IN2(n2660), .IN3(N18), .QN(n2659) );
  AO21X1 U2690 ( .IN1(N18), .IN2(N426), .IN3(n2660), .Q(n2603) );
  NAND2X0 U2691 ( .IN1(n2604), .IN2(n2661), .QN(n2660) );
  NAND3X0 U2692 ( .IN1(n2662), .IN2(n2663), .IN3(n2664), .QN(n2661) );
  AO21X1 U2693 ( .IN1(n2662), .IN2(n2663), .IN3(n2664), .Q(n2604) );
  NAND2X0 U2694 ( .IN1(n2609), .IN2(n2665), .QN(n2664) );
  NAND3X0 U2695 ( .IN1(N409), .IN2(n2666), .IN3(N35), .QN(n2665) );
  AO21X1 U2696 ( .IN1(N35), .IN2(N409), .IN3(n2666), .Q(n2609) );
  NAND2X0 U2697 ( .IN1(n2610), .IN2(n2667), .QN(n2666) );
  NAND3X0 U2698 ( .IN1(n2668), .IN2(n2669), .IN3(n2670), .QN(n2667) );
  AO21X1 U2699 ( .IN1(n2668), .IN2(n2669), .IN3(n2670), .Q(n2610) );
  NAND2X0 U2700 ( .IN1(n2615), .IN2(n2671), .QN(n2670) );
  NAND3X0 U2701 ( .IN1(N392), .IN2(n2672), .IN3(N52), .QN(n2671) );
  AO21X1 U2702 ( .IN1(N52), .IN2(N392), .IN3(n2672), .Q(n2615) );
  NAND2X0 U2703 ( .IN1(n2616), .IN2(n2673), .QN(n2672) );
  NAND3X0 U2704 ( .IN1(n2674), .IN2(n2675), .IN3(n2676), .QN(n2673) );
  AO21X1 U2705 ( .IN1(n2674), .IN2(n2675), .IN3(n2676), .Q(n2616) );
  XNOR2X1 U2706 ( .IN1(n2677), .IN2(keyinput15), .Q(n2676) );
  NAND2X0 U2707 ( .IN1(n2621), .IN2(n2678), .QN(n2677) );
  NAND3X0 U2708 ( .IN1(N375), .IN2(n2679), .IN3(N69), .QN(n2678) );
  AO21X1 U2709 ( .IN1(N69), .IN2(N375), .IN3(n2679), .Q(n2621) );
  NAND2X0 U2710 ( .IN1(n2622), .IN2(n2680), .QN(n2679) );
  NAND3X0 U2711 ( .IN1(n2681), .IN2(n2682), .IN3(n2683), .QN(n2680) );
  AO21X1 U2712 ( .IN1(n2681), .IN2(n2682), .IN3(n2683), .Q(n2622) );
  NAND2X0 U2713 ( .IN1(n2627), .IN2(n2684), .QN(n2683) );
  NAND3X0 U2714 ( .IN1(N358), .IN2(n2685), .IN3(N86), .QN(n2684) );
  AO21X1 U2715 ( .IN1(N86), .IN2(N358), .IN3(n2685), .Q(n2627) );
  NAND2X0 U2716 ( .IN1(n2628), .IN2(n2686), .QN(n2685) );
  NAND3X0 U2717 ( .IN1(n2687), .IN2(n2688), .IN3(n2689), .QN(n2686) );
  AO21X1 U2718 ( .IN1(n2687), .IN2(n2688), .IN3(n2689), .Q(n2628) );
  NAND2X0 U2719 ( .IN1(n2633), .IN2(n2690), .QN(n2689) );
  NAND3X0 U2720 ( .IN1(N341), .IN2(n2691), .IN3(N103), .QN(n2690) );
  AO21X1 U2721 ( .IN1(N103), .IN2(N341), .IN3(n2691), .Q(n2633) );
  NAND2X0 U2722 ( .IN1(n2634), .IN2(n2692), .QN(n2691) );
  NAND3X0 U2723 ( .IN1(n2693), .IN2(n2694), .IN3(n2695), .QN(n2692) );
  AO21X1 U2724 ( .IN1(n2693), .IN2(n2694), .IN3(n2695), .Q(n2634) );
  NAND2X0 U2725 ( .IN1(n2639), .IN2(n2696), .QN(n2695) );
  NAND3X0 U2726 ( .IN1(N324), .IN2(n2697), .IN3(N120), .QN(n2696) );
  AO21X1 U2727 ( .IN1(N120), .IN2(N324), .IN3(n2697), .Q(n2639) );
  NAND2X0 U2728 ( .IN1(n2640), .IN2(n2698), .QN(n2697) );
  NAND3X0 U2729 ( .IN1(n2699), .IN2(n2700), .IN3(n2701), .QN(n2698) );
  AO21X1 U2730 ( .IN1(n2699), .IN2(n2700), .IN3(n2701), .Q(n2640) );
  NAND2X0 U2731 ( .IN1(n2645), .IN2(n2702), .QN(n2701) );
  NAND3X0 U2732 ( .IN1(N307), .IN2(n2703), .IN3(N137), .QN(n2702) );
  AO21X1 U2733 ( .IN1(N137), .IN2(N307), .IN3(n2703), .Q(n2645) );
  OAI21X1 U2734 ( .IN1(n2704), .IN2(n2652), .IN3(n2646), .QN(n2703) );
  AO21X1 U2735 ( .IN1(n2705), .IN2(n2650), .IN3(n2706), .Q(n2646) );
  AO22X1 U2736 ( .IN1(N154), .IN2(N290), .IN3(N171), .IN4(N273), .Q(n2705) );
  INVX0 U2737 ( .INP(n2650), .ZN(n2652) );
  NAND3X0 U2738 ( .IN1(N171), .IN2(n2364), .IN3(N154), .QN(n2650) );
  NAND2X0 U2739 ( .IN1(n2656), .IN2(n2707), .QN(N4241) );
  NAND3X0 U2740 ( .IN1(N426), .IN2(n2708), .IN3(N1), .QN(n2707) );
  AO21X1 U2741 ( .IN1(N1), .IN2(N426), .IN3(n2708), .Q(n2656) );
  NAND2X0 U2742 ( .IN1(n2657), .IN2(n2709), .QN(n2708) );
  NAND3X0 U2743 ( .IN1(n2710), .IN2(n2711), .IN3(n2712), .QN(n2709) );
  AO21X1 U2744 ( .IN1(n2710), .IN2(n2711), .IN3(n2712), .Q(n2657) );
  NAND2X0 U2745 ( .IN1(n2662), .IN2(n2713), .QN(n2712) );
  NAND3X0 U2746 ( .IN1(N409), .IN2(n2714), .IN3(N18), .QN(n2713) );
  AO21X1 U2747 ( .IN1(N18), .IN2(N409), .IN3(n2714), .Q(n2662) );
  NAND2X0 U2748 ( .IN1(n2663), .IN2(n2715), .QN(n2714) );
  NAND3X0 U2749 ( .IN1(n2716), .IN2(n2717), .IN3(n2718), .QN(n2715) );
  AO21X1 U2750 ( .IN1(n2716), .IN2(n2717), .IN3(n2718), .Q(n2663) );
  NAND2X0 U2751 ( .IN1(n2668), .IN2(n2719), .QN(n2718) );
  NAND3X0 U2752 ( .IN1(N392), .IN2(n2720), .IN3(N35), .QN(n2719) );
  AO21X1 U2753 ( .IN1(N35), .IN2(N392), .IN3(n2720), .Q(n2668) );
  NAND2X0 U2754 ( .IN1(n2669), .IN2(n2721), .QN(n2720) );
  NAND3X0 U2755 ( .IN1(n2722), .IN2(n2723), .IN3(n2724), .QN(n2721) );
  AO21X1 U2756 ( .IN1(n2722), .IN2(n2723), .IN3(n2724), .Q(n2669) );
  NAND2X0 U2757 ( .IN1(n2674), .IN2(n2725), .QN(n2724) );
  NAND3X0 U2758 ( .IN1(N375), .IN2(n2726), .IN3(N52), .QN(n2725) );
  AO21X1 U2759 ( .IN1(N52), .IN2(N375), .IN3(n2726), .Q(n2674) );
  NAND2X0 U2760 ( .IN1(n2675), .IN2(n2727), .QN(n2726) );
  NAND3X0 U2761 ( .IN1(n2728), .IN2(n2729), .IN3(n2730), .QN(n2727) );
  AO21X1 U2762 ( .IN1(n2730), .IN2(n2729), .IN3(n2728), .Q(n2675) );
  NAND2X0 U2763 ( .IN1(n2681), .IN2(n2731), .QN(n2728) );
  NAND3X0 U2764 ( .IN1(N358), .IN2(n2732), .IN3(N69), .QN(n2731) );
  AO21X1 U2765 ( .IN1(N69), .IN2(N358), .IN3(n2732), .Q(n2681) );
  NAND2X0 U2766 ( .IN1(n2682), .IN2(n2733), .QN(n2732) );
  NAND3X0 U2767 ( .IN1(n2734), .IN2(n2735), .IN3(n2736), .QN(n2733) );
  AO21X1 U2768 ( .IN1(n2734), .IN2(n2735), .IN3(n2736), .Q(n2682) );
  NAND2X0 U2769 ( .IN1(n2687), .IN2(n2737), .QN(n2736) );
  NAND3X0 U2770 ( .IN1(N341), .IN2(n2738), .IN3(N86), .QN(n2737) );
  AO21X1 U2771 ( .IN1(N86), .IN2(N341), .IN3(n2738), .Q(n2687) );
  NAND2X0 U2772 ( .IN1(n2688), .IN2(n2739), .QN(n2738) );
  NAND3X0 U2773 ( .IN1(n2740), .IN2(n2741), .IN3(n2742), .QN(n2739) );
  AO21X1 U2774 ( .IN1(n2740), .IN2(n2741), .IN3(n2742), .Q(n2688) );
  NAND2X0 U2775 ( .IN1(n2693), .IN2(n2743), .QN(n2742) );
  NAND3X0 U2776 ( .IN1(N324), .IN2(n2744), .IN3(N103), .QN(n2743) );
  AO21X1 U2777 ( .IN1(N103), .IN2(N324), .IN3(n2744), .Q(n2693) );
  NAND2X0 U2778 ( .IN1(n2694), .IN2(n2745), .QN(n2744) );
  NAND3X0 U2779 ( .IN1(n2746), .IN2(n2747), .IN3(n2748), .QN(n2745) );
  AO21X1 U2780 ( .IN1(n2746), .IN2(n2747), .IN3(n2748), .Q(n2694) );
  NAND2X0 U2781 ( .IN1(n2699), .IN2(n2749), .QN(n2748) );
  NAND3X0 U2782 ( .IN1(N307), .IN2(n2750), .IN3(N120), .QN(n2749) );
  AO21X1 U2783 ( .IN1(N120), .IN2(N307), .IN3(n2750), .Q(n2699) );
  OAI21X1 U2784 ( .IN1(n2751), .IN2(n2706), .IN3(n2700), .QN(n2750) );
  AO21X1 U2785 ( .IN1(n2752), .IN2(n2704), .IN3(n2753), .Q(n2700) );
  AO22X1 U2786 ( .IN1(N137), .IN2(N290), .IN3(N154), .IN4(N273), .Q(n2752) );
  INVX0 U2787 ( .INP(n2704), .ZN(n2706) );
  NAND3X0 U2788 ( .IN1(N154), .IN2(n2364), .IN3(N137), .QN(n2704) );
  NAND2X0 U2789 ( .IN1(n2710), .IN2(n2754), .QN(N3895) );
  NAND3X0 U2790 ( .IN1(N409), .IN2(n2755), .IN3(N1), .QN(n2754) );
  AO21X1 U2791 ( .IN1(N1), .IN2(N409), .IN3(n2755), .Q(n2710) );
  NAND2X0 U2792 ( .IN1(n2711), .IN2(n2756), .QN(n2755) );
  NAND3X0 U2793 ( .IN1(n2757), .IN2(n2758), .IN3(n2759), .QN(n2756) );
  AO21X1 U2794 ( .IN1(n2757), .IN2(n2758), .IN3(n2759), .Q(n2711) );
  NAND2X0 U2795 ( .IN1(n2716), .IN2(n2760), .QN(n2759) );
  NAND3X0 U2796 ( .IN1(N392), .IN2(n2761), .IN3(N18), .QN(n2760) );
  AO21X1 U2797 ( .IN1(N18), .IN2(N392), .IN3(n2761), .Q(n2716) );
  NAND2X0 U2798 ( .IN1(n2717), .IN2(n2762), .QN(n2761) );
  NAND3X0 U2799 ( .IN1(n2763), .IN2(n2764), .IN3(n2765), .QN(n2762) );
  AO21X1 U2800 ( .IN1(n2763), .IN2(n2764), .IN3(n2765), .Q(n2717) );
  NAND2X0 U2801 ( .IN1(n2722), .IN2(n2766), .QN(n2765) );
  NAND3X0 U2802 ( .IN1(N375), .IN2(n2767), .IN3(N35), .QN(n2766) );
  AO21X1 U2803 ( .IN1(N35), .IN2(N375), .IN3(n2767), .Q(n2722) );
  NAND2X0 U2804 ( .IN1(n2723), .IN2(n2768), .QN(n2767) );
  NAND3X0 U2805 ( .IN1(n2769), .IN2(n2770), .IN3(n2771), .QN(n2768) );
  AO21X1 U2806 ( .IN1(n2769), .IN2(n2770), .IN3(n2771), .Q(n2723) );
  NAND2X0 U2807 ( .IN1(n2729), .IN2(n2772), .QN(n2771) );
  NAND3X0 U2808 ( .IN1(N358), .IN2(n2773), .IN3(N52), .QN(n2772) );
  AO21X1 U2809 ( .IN1(N52), .IN2(N358), .IN3(n2773), .Q(n2729) );
  NAND2X0 U2810 ( .IN1(n2730), .IN2(n2774), .QN(n2773) );
  NAND3X0 U2811 ( .IN1(n2775), .IN2(n2776), .IN3(n2777), .QN(n2774) );
  XOR2X1 U2812 ( .IN1(keyinput10), .IN2(n2778), .Q(n2730) );
  AOI21X1 U2813 ( .IN1(n2776), .IN2(n2775), .IN3(n2777), .QN(n2778) );
  NAND2X0 U2814 ( .IN1(n2734), .IN2(n2779), .QN(n2777) );
  NAND3X0 U2815 ( .IN1(N341), .IN2(n2780), .IN3(N69), .QN(n2779) );
  AO21X1 U2816 ( .IN1(N69), .IN2(N341), .IN3(n2780), .Q(n2734) );
  NAND2X0 U2817 ( .IN1(n2735), .IN2(n2781), .QN(n2780) );
  NAND3X0 U2818 ( .IN1(n2782), .IN2(n2783), .IN3(n2784), .QN(n2781) );
  AO21X1 U2819 ( .IN1(n2782), .IN2(n2783), .IN3(n2784), .Q(n2735) );
  NAND2X0 U2820 ( .IN1(n2740), .IN2(n2785), .QN(n2784) );
  NAND3X0 U2821 ( .IN1(N324), .IN2(n2786), .IN3(N86), .QN(n2785) );
  AO21X1 U2822 ( .IN1(N86), .IN2(N324), .IN3(n2786), .Q(n2740) );
  NAND2X0 U2823 ( .IN1(n2741), .IN2(n2787), .QN(n2786) );
  NAND3X0 U2824 ( .IN1(n2788), .IN2(n2789), .IN3(n2790), .QN(n2787) );
  AO21X1 U2825 ( .IN1(n2788), .IN2(n2789), .IN3(n2790), .Q(n2741) );
  NAND2X0 U2826 ( .IN1(n2746), .IN2(n2791), .QN(n2790) );
  NAND3X0 U2827 ( .IN1(N307), .IN2(n2792), .IN3(N103), .QN(n2791) );
  AO21X1 U2828 ( .IN1(N103), .IN2(N307), .IN3(n2792), .Q(n2746) );
  OAI21X1 U2829 ( .IN1(n2793), .IN2(n2753), .IN3(n2747), .QN(n2792) );
  AO21X1 U2830 ( .IN1(n2794), .IN2(n2751), .IN3(n2795), .Q(n2747) );
  AO22X1 U2831 ( .IN1(N120), .IN2(N290), .IN3(N137), .IN4(N273), .Q(n2794) );
  INVX0 U2832 ( .INP(n2751), .ZN(n2753) );
  NAND3X0 U2833 ( .IN1(N137), .IN2(n2364), .IN3(N120), .QN(n2751) );
  NAND2X0 U2834 ( .IN1(n2757), .IN2(n2796), .QN(N3552) );
  NAND3X0 U2835 ( .IN1(N392), .IN2(n2797), .IN3(N1), .QN(n2796) );
  AO21X1 U2836 ( .IN1(N1), .IN2(N392), .IN3(n2797), .Q(n2757) );
  NAND2X0 U2837 ( .IN1(n2758), .IN2(n2798), .QN(n2797) );
  NAND3X0 U2838 ( .IN1(n2799), .IN2(n2800), .IN3(n2801), .QN(n2798) );
  AO21X1 U2839 ( .IN1(n2799), .IN2(n2800), .IN3(n2801), .Q(n2758) );
  NAND2X0 U2840 ( .IN1(n2763), .IN2(n2802), .QN(n2801) );
  NAND3X0 U2841 ( .IN1(N375), .IN2(n2803), .IN3(N18), .QN(n2802) );
  AO21X1 U2842 ( .IN1(N18), .IN2(N375), .IN3(n2803), .Q(n2763) );
  NAND2X0 U2843 ( .IN1(n2764), .IN2(n2804), .QN(n2803) );
  NAND3X0 U2844 ( .IN1(n2805), .IN2(n2806), .IN3(n2807), .QN(n2804) );
  AO21X1 U2845 ( .IN1(n2805), .IN2(n2806), .IN3(n2807), .Q(n2764) );
  NAND2X0 U2846 ( .IN1(n2769), .IN2(n2808), .QN(n2807) );
  NAND3X0 U2847 ( .IN1(N358), .IN2(n2809), .IN3(N35), .QN(n2808) );
  AO21X1 U2848 ( .IN1(N35), .IN2(N358), .IN3(n2809), .Q(n2769) );
  NAND2X0 U2849 ( .IN1(n2770), .IN2(n2810), .QN(n2809) );
  NAND3X0 U2850 ( .IN1(n2811), .IN2(n2812), .IN3(n2813), .QN(n2810) );
  AO21X1 U2851 ( .IN1(n2811), .IN2(n2812), .IN3(n2813), .Q(n2770) );
  NAND2X0 U2852 ( .IN1(n2775), .IN2(n2814), .QN(n2813) );
  NAND3X0 U2853 ( .IN1(N341), .IN2(n2815), .IN3(N52), .QN(n2814) );
  AO21X1 U2854 ( .IN1(N52), .IN2(N341), .IN3(n2815), .Q(n2775) );
  NAND2X0 U2855 ( .IN1(n2776), .IN2(n2816), .QN(n2815) );
  NAND3X0 U2856 ( .IN1(n2817), .IN2(n2818), .IN3(n2819), .QN(n2816) );
  AO21X1 U2857 ( .IN1(n2819), .IN2(n2818), .IN3(n2817), .Q(n2776) );
  NAND2X0 U2858 ( .IN1(n2782), .IN2(n2820), .QN(n2817) );
  NAND3X0 U2859 ( .IN1(N324), .IN2(n2821), .IN3(N69), .QN(n2820) );
  AO21X1 U2860 ( .IN1(N69), .IN2(N324), .IN3(n2821), .Q(n2782) );
  NAND2X0 U2861 ( .IN1(n2783), .IN2(n2822), .QN(n2821) );
  NAND3X0 U2862 ( .IN1(n2823), .IN2(n2824), .IN3(n2825), .QN(n2822) );
  AO21X1 U2863 ( .IN1(n2823), .IN2(n2824), .IN3(n2825), .Q(n2783) );
  NAND2X0 U2864 ( .IN1(n2788), .IN2(n2826), .QN(n2825) );
  NAND3X0 U2865 ( .IN1(N307), .IN2(n2827), .IN3(N86), .QN(n2826) );
  AO21X1 U2866 ( .IN1(N86), .IN2(N307), .IN3(n2827), .Q(n2788) );
  OAI21X1 U2867 ( .IN1(n2828), .IN2(n2795), .IN3(n2789), .QN(n2827) );
  AO21X1 U2868 ( .IN1(n2829), .IN2(n2793), .IN3(n2830), .Q(n2789) );
  INVX0 U2869 ( .INP(n2828), .ZN(n2830) );
  AO22X1 U2870 ( .IN1(N103), .IN2(N290), .IN3(N120), .IN4(N273), .Q(n2829) );
  INVX0 U2871 ( .INP(n2793), .ZN(n2795) );
  NAND3X0 U2872 ( .IN1(N120), .IN2(n2364), .IN3(N103), .QN(n2793) );
  INVX0 U2873 ( .INP(n2831), .ZN(n2800) );
  NAND2X0 U2874 ( .IN1(n2799), .IN2(n2832), .QN(N3211) );
  NAND3X0 U2875 ( .IN1(N375), .IN2(n2833), .IN3(N1), .QN(n2832) );
  AO21X1 U2876 ( .IN1(N1), .IN2(N375), .IN3(n2833), .Q(n2799) );
  AO21X1 U2877 ( .IN1(n2834), .IN2(n2835), .IN3(n2831), .Q(n2833) );
  NOR2X0 U2878 ( .IN1(n2834), .IN2(n2835), .QN(n2831) );
  NAND2X0 U2879 ( .IN1(n2805), .IN2(n2836), .QN(n2835) );
  NAND3X0 U2880 ( .IN1(N358), .IN2(n2837), .IN3(N18), .QN(n2836) );
  AO21X1 U2881 ( .IN1(N18), .IN2(N358), .IN3(n2837), .Q(n2805) );
  NAND2X0 U2882 ( .IN1(n2806), .IN2(n2838), .QN(n2837) );
  NAND3X0 U2883 ( .IN1(n2839), .IN2(n2840), .IN3(n2841), .QN(n2838) );
  AO21X1 U2884 ( .IN1(n2839), .IN2(n2840), .IN3(n2841), .Q(n2806) );
  NAND2X0 U2885 ( .IN1(n2811), .IN2(n2842), .QN(n2841) );
  NAND3X0 U2886 ( .IN1(N341), .IN2(n2843), .IN3(N35), .QN(n2842) );
  AO21X1 U2887 ( .IN1(N35), .IN2(N341), .IN3(n2843), .Q(n2811) );
  NAND2X0 U2888 ( .IN1(n2812), .IN2(n2844), .QN(n2843) );
  NAND3X0 U2889 ( .IN1(n2845), .IN2(n2846), .IN3(n2847), .QN(n2844) );
  AO21X1 U2890 ( .IN1(n2845), .IN2(n2846), .IN3(n2847), .Q(n2812) );
  NAND2X0 U2891 ( .IN1(n2818), .IN2(n2848), .QN(n2847) );
  NAND3X0 U2892 ( .IN1(N324), .IN2(n2849), .IN3(N52), .QN(n2848) );
  AO21X1 U2893 ( .IN1(N52), .IN2(N324), .IN3(n2849), .Q(n2818) );
  AO21X1 U2894 ( .IN1(n2850), .IN2(n2851), .IN3(n2852), .Q(n2849) );
  INVX0 U2895 ( .INP(n2819), .ZN(n2852) );
  XNOR2X1 U2896 ( .IN1(n2853), .IN2(keyinput9), .Q(n2819) );
  OR2X1 U2897 ( .IN1(n2851), .IN2(n2850), .Q(n2853) );
  NAND2X0 U2898 ( .IN1(n2823), .IN2(n2854), .QN(n2851) );
  NAND3X0 U2899 ( .IN1(N307), .IN2(n2855), .IN3(N69), .QN(n2854) );
  AO21X1 U2900 ( .IN1(N69), .IN2(N307), .IN3(n2855), .Q(n2823) );
  AO21X1 U2901 ( .IN1(n2856), .IN2(n2857), .IN3(n2858), .Q(n2855) );
  INVX0 U2902 ( .INP(n2824), .ZN(n2858) );
  NAND2X0 U2903 ( .IN1(n2859), .IN2(n2860), .QN(n2824) );
  XOR2X1 U2904 ( .IN1(n2861), .IN2(keyinput4), .Q(n2859) );
  XNOR2X1 U2905 ( .IN1(keyinput4), .IN2(n2861), .Q(n2857) );
  NAND2X0 U2906 ( .IN1(n2862), .IN2(n2828), .QN(n2861) );
  NAND3X0 U2907 ( .IN1(N103), .IN2(n2364), .IN3(N86), .QN(n2828) );
  AO22X1 U2908 ( .IN1(N86), .IN2(N290), .IN3(N103), .IN4(N273), .Q(n2862) );
  AND2X1 U2909 ( .IN1(n2863), .IN2(n2864), .Q(n2850) );
  XOR2X1 U2910 ( .IN1(n2865), .IN2(keyinput11), .Q(n2834) );
  OA21X1 U2911 ( .IN1(n2866), .IN2(n2867), .IN3(n2868), .Q(n2865) );
  NAND2X0 U2912 ( .IN1(n2868), .IN2(n2869), .QN(N2877) );
  NAND3X0 U2913 ( .IN1(N358), .IN2(n2870), .IN3(N1), .QN(n2869) );
  AO21X1 U2914 ( .IN1(N1), .IN2(N358), .IN3(n2870), .Q(n2868) );
  XNOR2X1 U2915 ( .IN1(n2866), .IN2(n2867), .Q(n2870) );
  AND2X1 U2916 ( .IN1(n2871), .IN2(n2872), .Q(n2867) );
  NAND2X0 U2917 ( .IN1(n2839), .IN2(n2873), .QN(n2866) );
  NAND3X0 U2918 ( .IN1(N341), .IN2(n2874), .IN3(N18), .QN(n2873) );
  AO21X1 U2919 ( .IN1(N18), .IN2(N341), .IN3(n2874), .Q(n2839) );
  NAND2X0 U2920 ( .IN1(n2840), .IN2(n2875), .QN(n2874) );
  NAND3X0 U2921 ( .IN1(n2876), .IN2(n2877), .IN3(n2878), .QN(n2875) );
  AO21X1 U2922 ( .IN1(n2876), .IN2(n2877), .IN3(n2878), .Q(n2840) );
  NAND2X0 U2923 ( .IN1(n2845), .IN2(n2879), .QN(n2878) );
  NAND3X0 U2924 ( .IN1(N324), .IN2(n2880), .IN3(N35), .QN(n2879) );
  AO21X1 U2925 ( .IN1(N35), .IN2(N324), .IN3(n2880), .Q(n2845) );
  NAND2X0 U2926 ( .IN1(n2846), .IN2(n2881), .QN(n2880) );
  NAND3X0 U2927 ( .IN1(n2882), .IN2(n2883), .IN3(n2884), .QN(n2881) );
  AO21X1 U2928 ( .IN1(n2882), .IN2(n2883), .IN3(n2884), .Q(n2846) );
  NAND2X0 U2929 ( .IN1(n2863), .IN2(n2885), .QN(n2884) );
  NAND3X0 U2930 ( .IN1(N307), .IN2(n2886), .IN3(N52), .QN(n2885) );
  XNOR2X1 U2931 ( .IN1(keyinput6), .IN2(n2887), .Q(n2863) );
  AO21X1 U2932 ( .IN1(N52), .IN2(N307), .IN3(n2886), .Q(n2887) );
  OAI21X1 U2933 ( .IN1(n2888), .IN2(n2856), .IN3(n2864), .QN(n2886) );
  NAND2X0 U2934 ( .IN1(n2889), .IN2(n2888), .QN(n2864) );
  AO221X1 U2935 ( .IN1(n2890), .IN2(n2451), .IN3(n2890), .IN4(n2891), .IN5(
        n2856), .Q(n2889) );
  INVX0 U2936 ( .INP(N86), .ZN(n2891) );
  NAND2X0 U2937 ( .IN1(N69), .IN2(N290), .QN(n2890) );
  INVX0 U2938 ( .INP(n2860), .ZN(n2856) );
  NAND3X0 U2939 ( .IN1(N86), .IN2(n2364), .IN3(N69), .QN(n2860) );
  NAND2X0 U2940 ( .IN1(n2872), .IN2(n2892), .QN(N2548) );
  NAND3X0 U2941 ( .IN1(N341), .IN2(n2893), .IN3(N1), .QN(n2892) );
  AO21X1 U2942 ( .IN1(N1), .IN2(N341), .IN3(n2893), .Q(n2872) );
  NAND2X0 U2943 ( .IN1(n2871), .IN2(n2894), .QN(n2893) );
  NAND3X0 U2944 ( .IN1(n2895), .IN2(n2896), .IN3(n2897), .QN(n2894) );
  AO21X1 U2945 ( .IN1(n2895), .IN2(n2896), .IN3(n2897), .Q(n2871) );
  NAND2X0 U2946 ( .IN1(n2876), .IN2(n2898), .QN(n2897) );
  NAND3X0 U2947 ( .IN1(N324), .IN2(n2899), .IN3(N18), .QN(n2898) );
  AO21X1 U2948 ( .IN1(N18), .IN2(N324), .IN3(n2899), .Q(n2876) );
  NAND2X0 U2949 ( .IN1(n2877), .IN2(n2900), .QN(n2899) );
  NAND3X0 U2950 ( .IN1(n2901), .IN2(n2902), .IN3(n2903), .QN(n2900) );
  AO21X1 U2951 ( .IN1(n2901), .IN2(n2902), .IN3(n2903), .Q(n2877) );
  NAND2X0 U2952 ( .IN1(n2882), .IN2(n2904), .QN(n2903) );
  NAND3X0 U2953 ( .IN1(N307), .IN2(n2905), .IN3(N35), .QN(n2904) );
  AO21X1 U2954 ( .IN1(N35), .IN2(N307), .IN3(n2905), .Q(n2882) );
  AO21X1 U2955 ( .IN1(n2906), .IN2(n2888), .IN3(n2907), .Q(n2905) );
  INVX0 U2956 ( .INP(n2883), .ZN(n2907) );
  AO21X1 U2957 ( .IN1(n2908), .IN2(n2888), .IN3(n2906), .Q(n2883) );
  AO22X1 U2958 ( .IN1(N52), .IN2(N290), .IN3(N69), .IN4(N273), .Q(n2908) );
  NAND3X0 U2959 ( .IN1(N69), .IN2(n2364), .IN3(N52), .QN(n2888) );
  NAND2X0 U2960 ( .IN1(n2895), .IN2(n2909), .QN(N2223) );
  NAND3X0 U2961 ( .IN1(N324), .IN2(n2910), .IN3(N1), .QN(n2909) );
  AO21X1 U2962 ( .IN1(N1), .IN2(N324), .IN3(n2910), .Q(n2895) );
  NAND2X0 U2963 ( .IN1(n2896), .IN2(n2911), .QN(n2910) );
  NAND3X0 U2964 ( .IN1(n2912), .IN2(n2913), .IN3(n2914), .QN(n2911) );
  AO21X1 U2965 ( .IN1(n2912), .IN2(n2913), .IN3(n2914), .Q(n2896) );
  NAND2X0 U2966 ( .IN1(n2901), .IN2(n2915), .QN(n2914) );
  NAND3X0 U2967 ( .IN1(N307), .IN2(n2916), .IN3(N18), .QN(n2915) );
  AO21X1 U2968 ( .IN1(N18), .IN2(N307), .IN3(n2916), .Q(n2901) );
  OAI21X1 U2969 ( .IN1(n2917), .IN2(n2906), .IN3(n2902), .QN(n2916) );
  AO21X1 U2970 ( .IN1(n2918), .IN2(n2919), .IN3(n2920), .Q(n2902) );
  INVX0 U2971 ( .INP(n2917), .ZN(n2920) );
  AO22X1 U2972 ( .IN1(N35), .IN2(N290), .IN3(N52), .IN4(N273), .Q(n2918) );
  INVX0 U2973 ( .INP(n2919), .ZN(n2906) );
  NAND3X0 U2974 ( .IN1(N52), .IN2(n2364), .IN3(N35), .QN(n2919) );
  NAND2X0 U2975 ( .IN1(n2912), .IN2(n2921), .QN(N1901) );
  NAND3X0 U2976 ( .IN1(N307), .IN2(n2922), .IN3(N1), .QN(n2921) );
  AO21X1 U2977 ( .IN1(N1), .IN2(N307), .IN3(n2922), .Q(n2912) );
  AO21X1 U2978 ( .IN1(n2923), .IN2(n2917), .IN3(n2924), .Q(n2922) );
  INVX0 U2979 ( .INP(n2913), .ZN(n2924) );
  AO21X1 U2980 ( .IN1(n2925), .IN2(n2917), .IN3(n2923), .Q(n2913) );
  AO22X1 U2981 ( .IN1(N18), .IN2(N290), .IN3(N35), .IN4(N273), .Q(n2925) );
  NAND3X0 U2982 ( .IN1(N35), .IN2(n2364), .IN3(N18), .QN(n2917) );
  NOR2X0 U2983 ( .IN1(n2451), .IN2(n2926), .QN(n2364) );
  NOR2X0 U2984 ( .IN1(n2923), .IN2(n2927), .QN(N1581) );
  AOI22X1 U2985 ( .IN1(N273), .IN2(N18), .IN3(N290), .IN4(N1), .QN(n2927) );
  AND3X1 U2986 ( .IN1(N18), .IN2(n2452), .IN3(N545), .Q(n2923) );
  AND2X1 U2987 ( .IN1(N1), .IN2(N273), .Q(N545) );
  INVX0 U2988 ( .INP(n2926), .ZN(n2452) );
  NOR2X0 U2989 ( .IN1(n2451), .IN2(N290), .QN(n2926) );
  INVX0 U2990 ( .INP(N273), .ZN(n2451) );
endmodule

