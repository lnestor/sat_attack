`timescale 1ns / 1ps
// Verilog
// c499
// Ninputs 41
// Noutputs 32
// NtotalGates 202
// XOR2 104
// AND2 40
// NOT1 40
// AND4 8
// OR4 2
// AND5 8

module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
                  N753,N754,N755,
        keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4,
        keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9,
        keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14,
        keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19,
        keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24,
        keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29,
        keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34,
        keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39,
        keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44,
        keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49,
        keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54,
        keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59,
        keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64,
        keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69,
        keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74,
        keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79,
        keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84,
        keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89,
        keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94,
        keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99,
        keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104,
        keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109,
        keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114,
        keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119,
        keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124,
        keyIn_0_125, keyIn_0_126, keyIn_0_127);

  input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4;
  input keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9;
  input keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14;
  input keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19;
  input keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24;
  input keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29;
  input keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34;
  input keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39;
  input keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44;
  input keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49;
  input keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54;
  input keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59;
  input keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64;
  input keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69;
  input keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74;
  input keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79;
  input keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84;
  input keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89;
  input keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94;
  input keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99;
  input keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104;
  input keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109;
  input keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114;
  input keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119;
  input keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124;
  input keyIn_0_125, keyIn_0_126, keyIn_0_127;

  wire [0:127] KeyWire_0;
  wire [0:59] KeyNOTWire_0;

input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;

output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;

wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723;

xor XOR2_1 (N250, N1, N5);
xor XOR2_2 (N251, N9, N13);
  xor XOR2_3 (KeyWire_0[0], N17, N21);
  xnor KeyGate_0_0(N252, keyIn_0_0, KeyWire_0[0]);
xor XOR2_4 (N253, N25, N29);
  xor XOR2_5 (KeyWire_0[1], N33, N37);
  xor KeyGate_0_1(KeyNOTWire_0[0], keyIn_0_1, KeyWire_0[1]);
  not KeyNOTGate_0_0(N254, KeyNOTWire_0[0]);
  xor XOR2_6 (KeyWire_0[2], N41, N45);
  xor KeyGate_0_2(N255, keyIn_0_2, KeyWire_0[2]);
  xor XOR2_7 (KeyWire_0[3], N49, N53);
  xor KeyGate_0_3(KeyNOTWire_0[1], keyIn_0_3, KeyWire_0[3]);
  not KeyNOTGate_0_1(N256, KeyNOTWire_0[1]);
  xor XOR2_8 (KeyWire_0[4], N57, N61);
  xnor KeyGate_0_4(N257, keyIn_0_4, KeyWire_0[4]);
xor XOR2_9 (N258, N65, N69);
xor XOR2_10 (N259, N73, N77);
  xor XOR2_11 (KeyWire_0[5], N81, N85);
  xnor KeyGate_0_5(N260, keyIn_0_5, KeyWire_0[5]);
  xor XOR2_12 (KeyWire_0[6], N89, N93);
  xor KeyGate_0_6(N261, keyIn_0_6, KeyWire_0[6]);
xor XOR2_13 (N262, N97, N101);
  xor XOR2_14 (KeyWire_0[7], N105, N109);
  xor KeyGate_0_7(KeyNOTWire_0[2], keyIn_0_7, KeyWire_0[7]);
  not KeyNOTGate_0_2(N263, KeyNOTWire_0[2]);
xor XOR2_15 (N264, N113, N117);
  xor XOR2_16 (KeyWire_0[8], N121, N125);
  xor KeyGate_0_8(N265, keyIn_0_8, KeyWire_0[8]);
  and AND2_17 (KeyWire_0[9], N129, N137);
  xor KeyGate_0_9(KeyNOTWire_0[3], keyIn_0_9, KeyWire_0[9]);
  not KeyNOTGate_0_3(N266, KeyNOTWire_0[3]);
  and AND2_18 (KeyWire_0[10], N130, N137);
  xnor KeyGate_0_10(N267, keyIn_0_10, KeyWire_0[10]);
  and AND2_19 (KeyWire_0[11], N131, N137);
  xor KeyGate_0_11(KeyNOTWire_0[4], keyIn_0_11, KeyWire_0[11]);
  not KeyNOTGate_0_4(N268, KeyNOTWire_0[4]);
  and AND2_20 (KeyWire_0[12], N132, N137);
  xor KeyGate_0_12(KeyNOTWire_0[5], keyIn_0_12, KeyWire_0[12]);
  not KeyNOTGate_0_5(N269, KeyNOTWire_0[5]);
  and AND2_21 (KeyWire_0[13], N133, N137);
  xnor KeyGate_0_13(KeyNOTWire_0[6], keyIn_0_13, KeyWire_0[13]);
  not KeyNOTGate_0_6(N270, KeyNOTWire_0[6]);
  and AND2_22 (KeyWire_0[14], N134, N137);
  xnor KeyGate_0_14(KeyNOTWire_0[7], keyIn_0_14, KeyWire_0[14]);
  not KeyNOTGate_0_7(N271, KeyNOTWire_0[7]);
and AND2_23 (N272, N135, N137);
  and AND2_24 (KeyWire_0[15], N136, N137);
  xnor KeyGate_0_15(N273, keyIn_0_15, KeyWire_0[15]);
xor XOR2_25 (N274, N1, N17);
  xor XOR2_26 (KeyWire_0[16], N33, N49);
  xnor KeyGate_0_16(KeyNOTWire_0[8], keyIn_0_16, KeyWire_0[16]);
  not KeyNOTGate_0_8(N275, KeyNOTWire_0[8]);
  xor XOR2_27 (KeyWire_0[17], N5, N21);
  xnor KeyGate_0_17(N276, keyIn_0_17, KeyWire_0[17]);
  xor XOR2_28 (KeyWire_0[18], N37, N53);
  xnor KeyGate_0_18(N277, keyIn_0_18, KeyWire_0[18]);
xor XOR2_29 (N278, N9, N25);
  xor XOR2_30 (KeyWire_0[19], N41, N57);
  xnor KeyGate_0_19(N279, keyIn_0_19, KeyWire_0[19]);
  xor XOR2_31 (KeyWire_0[20], N13, N29);
  xnor KeyGate_0_20(N280, keyIn_0_20, KeyWire_0[20]);
xor XOR2_32 (N281, N45, N61);
  xor XOR2_33 (KeyWire_0[21], N65, N81);
  xor KeyGate_0_21(KeyNOTWire_0[9], keyIn_0_21, KeyWire_0[21]);
  not KeyNOTGate_0_9(N282, KeyNOTWire_0[9]);
  xor XOR2_34 (KeyWire_0[22], N97, N113);
  xnor KeyGate_0_22(N283, keyIn_0_22, KeyWire_0[22]);
  xor XOR2_35 (KeyWire_0[23], N69, N85);
  xor KeyGate_0_23(KeyNOTWire_0[10], keyIn_0_23, KeyWire_0[23]);
  not KeyNOTGate_0_10(N284, KeyNOTWire_0[10]);
  xor XOR2_36 (KeyWire_0[24], N101, N117);
  xor KeyGate_0_24(N285, keyIn_0_24, KeyWire_0[24]);
xor XOR2_37 (N286, N73, N89);
xor XOR2_38 (N287, N105, N121);
xor XOR2_39 (N288, N77, N93);
xor XOR2_40 (N289, N109, N125);
xor XOR2_41 (N290, N250, N251);
  xor XOR2_42 (KeyWire_0[25], N252, N253);
  xor KeyGate_0_25(KeyNOTWire_0[11], keyIn_0_25, KeyWire_0[25]);
  not KeyNOTGate_0_11(N293, KeyNOTWire_0[11]);
  xor XOR2_43 (KeyWire_0[26], N254, N255);
  xnor KeyGate_0_26(N296, keyIn_0_26, KeyWire_0[26]);
  xor XOR2_44 (KeyWire_0[27], N256, N257);
  xor KeyGate_0_27(N299, keyIn_0_27, KeyWire_0[27]);
xor XOR2_45 (N302, N258, N259);
  xor XOR2_46 (KeyWire_0[28], N260, N261);
  xnor KeyGate_0_28(KeyNOTWire_0[12], keyIn_0_28, KeyWire_0[28]);
  not KeyNOTGate_0_12(N305, KeyNOTWire_0[12]);
xor XOR2_47 (N308, N262, N263);
xor XOR2_48 (N311, N264, N265);
xor XOR2_49 (N314, N274, N275);
xor XOR2_50 (N315, N276, N277);
  xor XOR2_51 (KeyWire_0[29], N278, N279);
  xor KeyGate_0_29(KeyNOTWire_0[13], keyIn_0_29, KeyWire_0[29]);
  not KeyNOTGate_0_13(N316, KeyNOTWire_0[13]);
  xor XOR2_52 (KeyWire_0[30], N280, N281);
  xnor KeyGate_0_30(KeyNOTWire_0[14], keyIn_0_30, KeyWire_0[30]);
  not KeyNOTGate_0_14(N317, KeyNOTWire_0[14]);
xor XOR2_53 (N318, N282, N283);
xor XOR2_54 (N319, N284, N285);
  xor XOR2_55 (KeyWire_0[31], N286, N287);
  xor KeyGate_0_31(N320, keyIn_0_31, KeyWire_0[31]);
  xor XOR2_56 (KeyWire_0[32], N288, N289);
  xor KeyGate_0_32(KeyNOTWire_0[15], keyIn_0_32, KeyWire_0[32]);
  not KeyNOTGate_0_15(N321, KeyNOTWire_0[15]);
xor XOR2_57 (N338, N290, N293);
  xor XOR2_58 (KeyWire_0[33], N296, N299);
  xnor KeyGate_0_33(N339, keyIn_0_33, KeyWire_0[33]);
xor XOR2_59 (N340, N290, N296);
xor XOR2_60 (N341, N293, N299);
  xor XOR2_61 (KeyWire_0[34], N302, N305);
  xnor KeyGate_0_34(KeyNOTWire_0[16], keyIn_0_34, KeyWire_0[34]);
  not KeyNOTGate_0_16(N342, KeyNOTWire_0[16]);
  xor XOR2_62 (KeyWire_0[35], N308, N311);
  xor KeyGate_0_35(N343, keyIn_0_35, KeyWire_0[35]);
xor XOR2_63 (N344, N302, N308);
xor XOR2_64 (N345, N305, N311);
  xor XOR2_65 (KeyWire_0[36], N266, N342);
  xor KeyGate_0_36(N346, keyIn_0_36, KeyWire_0[36]);
xor XOR2_66 (N347, N267, N343);
xor XOR2_67 (N348, N268, N344);
  xor XOR2_68 (KeyWire_0[37], N269, N345);
  xnor KeyGate_0_37(KeyNOTWire_0[17], keyIn_0_37, KeyWire_0[37]);
  not KeyNOTGate_0_17(N349, KeyNOTWire_0[17]);
  xor XOR2_69 (KeyWire_0[38], N270, N338);
  xor KeyGate_0_38(KeyNOTWire_0[18], keyIn_0_38, KeyWire_0[38]);
  not KeyNOTGate_0_18(N350, KeyNOTWire_0[18]);
  xor XOR2_70 (KeyWire_0[39], N271, N339);
  xor KeyGate_0_39(N351, keyIn_0_39, KeyWire_0[39]);
xor XOR2_71 (N352, N272, N340);
xor XOR2_72 (N353, N273, N341);
  xor XOR2_73 (KeyWire_0[40], N314, N346);
  xnor KeyGate_0_40(KeyNOTWire_0[19], keyIn_0_40, KeyWire_0[40]);
  not KeyNOTGate_0_19(N354, KeyNOTWire_0[19]);
xor XOR2_74 (N367, N315, N347);
xor XOR2_75 (N380, N316, N348);
  xor XOR2_76 (KeyWire_0[41], N317, N349);
  xnor KeyGate_0_41(KeyNOTWire_0[20], keyIn_0_41, KeyWire_0[41]);
  not KeyNOTGate_0_20(N393, KeyNOTWire_0[20]);
  xor XOR2_77 (KeyWire_0[42], N318, N350);
  xnor KeyGate_0_42(KeyNOTWire_0[21], keyIn_0_42, KeyWire_0[42]);
  not KeyNOTGate_0_21(N406, KeyNOTWire_0[21]);
  xor XOR2_78 (KeyWire_0[43], N319, N351);
  xor KeyGate_0_43(KeyNOTWire_0[22], keyIn_0_43, KeyWire_0[43]);
  not KeyNOTGate_0_22(N419, KeyNOTWire_0[22]);
  xor XOR2_79 (KeyWire_0[44], N320, N352);
  xor KeyGate_0_44(N432, keyIn_0_44, KeyWire_0[44]);
  xor XOR2_80 (KeyWire_0[45], N321, N353);
  xnor KeyGate_0_45(N445, keyIn_0_45, KeyWire_0[45]);
  not NOT1_81 (KeyWire_0[46], N354);
  xnor KeyGate_0_46(N554, keyIn_0_46, KeyWire_0[46]);
  not NOT1_82 (KeyWire_0[47], N367);
  xnor KeyGate_0_47(N555, keyIn_0_47, KeyWire_0[47]);
  not NOT1_83 (KeyWire_0[48], N380);
  xnor KeyGate_0_48(N556, keyIn_0_48, KeyWire_0[48]);
  not NOT1_84 (KeyWire_0[49], N354);
  xnor KeyGate_0_49(N557, keyIn_0_49, KeyWire_0[49]);
  not NOT1_85 (KeyWire_0[50], N367);
  xnor KeyGate_0_50(N558, keyIn_0_50, KeyWire_0[50]);
not NOT1_86 (N559, N393);
not NOT1_87 (N560, N354);
  not NOT1_88 (KeyWire_0[51], N380);
  xnor KeyGate_0_51(N561, keyIn_0_51, KeyWire_0[51]);
  not NOT1_89 (KeyWire_0[52], N393);
  xnor KeyGate_0_52(KeyNOTWire_0[23], keyIn_0_52, KeyWire_0[52]);
  not KeyNOTGate_0_23(N562, KeyNOTWire_0[23]);
not NOT1_90 (N563, N367);
not NOT1_91 (N564, N380);
not NOT1_92 (N565, N393);
  not NOT1_93 (KeyWire_0[53], N419);
  xor KeyGate_0_53(N566, keyIn_0_53, KeyWire_0[53]);
  not NOT1_94 (KeyWire_0[54], N445);
  xnor KeyGate_0_54(KeyNOTWire_0[24], keyIn_0_54, KeyWire_0[54]);
  not KeyNOTGate_0_24(N567, KeyNOTWire_0[24]);
  not NOT1_95 (KeyWire_0[55], N419);
  xnor KeyGate_0_55(N568, keyIn_0_55, KeyWire_0[55]);
not NOT1_96 (N569, N432);
  not NOT1_97 (KeyWire_0[56], N406);
  xor KeyGate_0_56(KeyNOTWire_0[25], keyIn_0_56, KeyWire_0[56]);
  not KeyNOTGate_0_25(N570, KeyNOTWire_0[25]);
not NOT1_98 (N571, N445);
  not NOT1_99 (KeyWire_0[57], N406);
  xnor KeyGate_0_57(N572, keyIn_0_57, KeyWire_0[57]);
  not NOT1_100 (KeyWire_0[58], N432);
  xor KeyGate_0_58(N573, keyIn_0_58, KeyWire_0[58]);
not NOT1_101 (N574, N406);
  not NOT1_102 (KeyWire_0[59], N419);
  xnor KeyGate_0_59(KeyNOTWire_0[26], keyIn_0_59, KeyWire_0[59]);
  not KeyNOTGate_0_26(N575, KeyNOTWire_0[26]);
  not NOT1_103 (KeyWire_0[60], N432);
  xor KeyGate_0_60(N576, keyIn_0_60, KeyWire_0[60]);
not NOT1_104 (N577, N406);
not NOT1_105 (N578, N419);
  not NOT1_106 (KeyWire_0[61], N445);
  xor KeyGate_0_61(KeyNOTWire_0[27], keyIn_0_61, KeyWire_0[61]);
  not KeyNOTGate_0_27(N579, KeyNOTWire_0[27]);
  not NOT1_107 (KeyWire_0[62], N406);
  xor KeyGate_0_62(KeyNOTWire_0[28], keyIn_0_62, KeyWire_0[62]);
  not KeyNOTGate_0_28(N580, KeyNOTWire_0[28]);
  not NOT1_108 (KeyWire_0[63], N432);
  xor KeyGate_0_63(KeyNOTWire_0[29], keyIn_0_63, KeyWire_0[63]);
  not KeyNOTGate_0_29(N581, KeyNOTWire_0[29]);
  not NOT1_109 (KeyWire_0[64], N445);
  xor KeyGate_0_64(KeyNOTWire_0[30], keyIn_0_64, KeyWire_0[64]);
  not KeyNOTGate_0_30(N582, KeyNOTWire_0[30]);
not NOT1_110 (N583, N419);
  not NOT1_111 (KeyWire_0[65], N432);
  xnor KeyGate_0_65(KeyNOTWire_0[31], keyIn_0_65, KeyWire_0[65]);
  not KeyNOTGate_0_31(N584, KeyNOTWire_0[31]);
  not NOT1_112 (KeyWire_0[66], N445);
  xor KeyGate_0_66(N585, keyIn_0_66, KeyWire_0[66]);
  not NOT1_113 (KeyWire_0[67], N367);
  xnor KeyGate_0_67(KeyNOTWire_0[32], keyIn_0_67, KeyWire_0[67]);
  not KeyNOTGate_0_32(N586, KeyNOTWire_0[32]);
  not NOT1_114 (KeyWire_0[68], N393);
  xor KeyGate_0_68(KeyNOTWire_0[33], keyIn_0_68, KeyWire_0[68]);
  not KeyNOTGate_0_33(N587, KeyNOTWire_0[33]);
  not NOT1_115 (KeyWire_0[69], N367);
  xor KeyGate_0_69(N588, keyIn_0_69, KeyWire_0[69]);
  not NOT1_116 (KeyWire_0[70], N380);
  xor KeyGate_0_70(N589, keyIn_0_70, KeyWire_0[70]);
not NOT1_117 (N590, N354);
not NOT1_118 (N591, N393);
not NOT1_119 (N592, N354);
  not NOT1_120 (KeyWire_0[71], N380);
  xnor KeyGate_0_71(N593, keyIn_0_71, KeyWire_0[71]);
  and AND4_121 (KeyWire_0[72], N554, N555, N556, N393);
  xnor KeyGate_0_72(KeyNOTWire_0[34], keyIn_0_72, KeyWire_0[72]);
  not KeyNOTGate_0_34(N594, KeyNOTWire_0[34]);
  and AND4_122 (KeyWire_0[73], N557, N558, N380, N559);
  xnor KeyGate_0_73(KeyNOTWire_0[35], keyIn_0_73, KeyWire_0[73]);
  not KeyNOTGate_0_35(N595, KeyNOTWire_0[35]);
  and AND4_123 (KeyWire_0[74], N560, N367, N561, N562);
  xor KeyGate_0_74(N596, keyIn_0_74, KeyWire_0[74]);
  and AND4_124 (KeyWire_0[75], N354, N563, N564, N565);
  xor KeyGate_0_75(KeyNOTWire_0[36], keyIn_0_75, KeyWire_0[75]);
  not KeyNOTGate_0_36(N597, KeyNOTWire_0[36]);
  and AND4_125 (KeyWire_0[76], N574, N575, N576, N445);
  xor KeyGate_0_76(KeyNOTWire_0[37], keyIn_0_76, KeyWire_0[76]);
  not KeyNOTGate_0_37(N598, KeyNOTWire_0[37]);
and AND4_126 (N599, N577, N578, N432, N579);
and AND4_127 (N600, N580, N419, N581, N582);
  and AND4_128 (KeyWire_0[77], N406, N583, N584, N585);
  xnor KeyGate_0_77(N601, keyIn_0_77, KeyWire_0[77]);
  or OR4_129 (KeyWire_0[78], N594, N595, N596, N597);
  xnor KeyGate_0_78(N602, keyIn_0_78, KeyWire_0[78]);
  or OR4_130 (KeyWire_0[79], N598, N599, N600, N601);
  xnor KeyGate_0_79(N607, keyIn_0_79, KeyWire_0[79]);
and AND5_131 (N620, N406, N566, N432, N567, N602);
  and AND5_132 (KeyWire_0[80], N406, N568, N569, N445, N602);
  xor KeyGate_0_80(N625, keyIn_0_80, KeyWire_0[80]);
and AND5_133 (N630, N570, N419, N432, N571, N602);
  and AND5_134 (KeyWire_0[81], N572, N419, N573, N445, N602);
  xor KeyGate_0_81(KeyNOTWire_0[38], keyIn_0_81, KeyWire_0[81]);
  not KeyNOTGate_0_38(N635, KeyNOTWire_0[38]);
  and AND5_135 (KeyWire_0[82], N354, N586, N380, N587, N607);
  xor KeyGate_0_82(KeyNOTWire_0[39], keyIn_0_82, KeyWire_0[82]);
  not KeyNOTGate_0_39(N640, KeyNOTWire_0[39]);
  and AND5_136 (KeyWire_0[83], N354, N588, N589, N393, N607);
  xor KeyGate_0_83(N645, keyIn_0_83, KeyWire_0[83]);
  and AND5_137 (KeyWire_0[84], N590, N367, N380, N591, N607);
  xnor KeyGate_0_84(N650, keyIn_0_84, KeyWire_0[84]);
  and AND5_138 (KeyWire_0[85], N592, N367, N593, N393, N607);
  xnor KeyGate_0_85(KeyNOTWire_0[40], keyIn_0_85, KeyWire_0[85]);
  not KeyNOTGate_0_40(N655, KeyNOTWire_0[40]);
and AND2_139 (N692, N354, N620);
  and AND2_140 (KeyWire_0[86], N367, N620);
  xor KeyGate_0_86(KeyNOTWire_0[41], keyIn_0_86, KeyWire_0[86]);
  not KeyNOTGate_0_41(N693, KeyNOTWire_0[41]);
  and AND2_141 (KeyWire_0[87], N380, N620);
  xnor KeyGate_0_87(KeyNOTWire_0[42], keyIn_0_87, KeyWire_0[87]);
  not KeyNOTGate_0_42(N694, KeyNOTWire_0[42]);
  and AND2_142 (KeyWire_0[88], N393, N620);
  xor KeyGate_0_88(N695, keyIn_0_88, KeyWire_0[88]);
and AND2_143 (N696, N354, N625);
and AND2_144 (N697, N367, N625);
and AND2_145 (N698, N380, N625);
and AND2_146 (N699, N393, N625);
  and AND2_147 (KeyWire_0[89], N354, N630);
  xnor KeyGate_0_89(N700, keyIn_0_89, KeyWire_0[89]);
  and AND2_148 (KeyWire_0[90], N367, N630);
  xnor KeyGate_0_90(N701, keyIn_0_90, KeyWire_0[90]);
  and AND2_149 (KeyWire_0[91], N380, N630);
  xnor KeyGate_0_91(N702, keyIn_0_91, KeyWire_0[91]);
and AND2_150 (N703, N393, N630);
  and AND2_151 (KeyWire_0[92], N354, N635);
  xor KeyGate_0_92(KeyNOTWire_0[43], keyIn_0_92, KeyWire_0[92]);
  not KeyNOTGate_0_43(N704, KeyNOTWire_0[43]);
  and AND2_152 (KeyWire_0[93], N367, N635);
  xor KeyGate_0_93(KeyNOTWire_0[44], keyIn_0_93, KeyWire_0[93]);
  not KeyNOTGate_0_44(N705, KeyNOTWire_0[44]);
  and AND2_153 (KeyWire_0[94], N380, N635);
  xor KeyGate_0_94(KeyNOTWire_0[45], keyIn_0_94, KeyWire_0[94]);
  not KeyNOTGate_0_45(N706, KeyNOTWire_0[45]);
  and AND2_154 (KeyWire_0[95], N393, N635);
  xor KeyGate_0_95(N707, keyIn_0_95, KeyWire_0[95]);
  and AND2_155 (KeyWire_0[96], N406, N640);
  xnor KeyGate_0_96(KeyNOTWire_0[46], keyIn_0_96, KeyWire_0[96]);
  not KeyNOTGate_0_46(N708, KeyNOTWire_0[46]);
  and AND2_156 (KeyWire_0[97], N419, N640);
  xnor KeyGate_0_97(N709, keyIn_0_97, KeyWire_0[97]);
  and AND2_157 (KeyWire_0[98], N432, N640);
  xor KeyGate_0_98(N710, keyIn_0_98, KeyWire_0[98]);
and AND2_158 (N711, N445, N640);
  and AND2_159 (KeyWire_0[99], N406, N645);
  xor KeyGate_0_99(KeyNOTWire_0[47], keyIn_0_99, KeyWire_0[99]);
  not KeyNOTGate_0_47(N712, KeyNOTWire_0[47]);
and AND2_160 (N713, N419, N645);
  and AND2_161 (KeyWire_0[100], N432, N645);
  xor KeyGate_0_100(KeyNOTWire_0[48], keyIn_0_100, KeyWire_0[100]);
  not KeyNOTGate_0_48(N714, KeyNOTWire_0[48]);
  and AND2_162 (KeyWire_0[101], N445, N645);
  xor KeyGate_0_101(N715, keyIn_0_101, KeyWire_0[101]);
  and AND2_163 (KeyWire_0[102], N406, N650);
  xor KeyGate_0_102(N716, keyIn_0_102, KeyWire_0[102]);
  and AND2_164 (KeyWire_0[103], N419, N650);
  xnor KeyGate_0_103(KeyNOTWire_0[49], keyIn_0_103, KeyWire_0[103]);
  not KeyNOTGate_0_49(N717, KeyNOTWire_0[49]);
  and AND2_165 (KeyWire_0[104], N432, N650);
  xnor KeyGate_0_104(N718, keyIn_0_104, KeyWire_0[104]);
and AND2_166 (N719, N445, N650);
  and AND2_167 (KeyWire_0[105], N406, N655);
  xnor KeyGate_0_105(N720, keyIn_0_105, KeyWire_0[105]);
  and AND2_168 (KeyWire_0[106], N419, N655);
  xnor KeyGate_0_106(N721, keyIn_0_106, KeyWire_0[106]);
and AND2_169 (N722, N432, N655);
and AND2_170 (N723, N445, N655);
  xor XOR2_171 (KeyWire_0[107], N1, N692);
  xnor KeyGate_0_107(KeyNOTWire_0[50], keyIn_0_107, KeyWire_0[107]);
  not KeyNOTGate_0_50(N724, KeyNOTWire_0[50]);
  xor XOR2_172 (KeyWire_0[108], N5, N693);
  xor KeyGate_0_108(KeyNOTWire_0[51], keyIn_0_108, KeyWire_0[108]);
  not KeyNOTGate_0_51(N725, KeyNOTWire_0[51]);
  xor XOR2_173 (KeyWire_0[109], N9, N694);
  xnor KeyGate_0_109(N726, keyIn_0_109, KeyWire_0[109]);
  xor XOR2_174 (KeyWire_0[110], N13, N695);
  xnor KeyGate_0_110(N727, keyIn_0_110, KeyWire_0[110]);
xor XOR2_175 (N728, N17, N696);
xor XOR2_176 (N729, N21, N697);
xor XOR2_177 (N730, N25, N698);
  xor XOR2_178 (KeyWire_0[111], N29, N699);
  xor KeyGate_0_111(KeyNOTWire_0[52], keyIn_0_111, KeyWire_0[111]);
  not KeyNOTGate_0_52(N731, KeyNOTWire_0[52]);
  xor XOR2_179 (KeyWire_0[112], N33, N700);
  xnor KeyGate_0_112(N732, keyIn_0_112, KeyWire_0[112]);
  xor XOR2_180 (KeyWire_0[113], N37, N701);
  xor KeyGate_0_113(N733, keyIn_0_113, KeyWire_0[113]);
xor XOR2_181 (N734, N41, N702);
  xor XOR2_182 (KeyWire_0[114], N45, N703);
  xor KeyGate_0_114(N735, keyIn_0_114, KeyWire_0[114]);
xor XOR2_183 (N736, N49, N704);
xor XOR2_184 (N737, N53, N705);
  xor XOR2_185 (KeyWire_0[115], N57, N706);
  xor KeyGate_0_115(KeyNOTWire_0[53], keyIn_0_115, KeyWire_0[115]);
  not KeyNOTGate_0_53(N738, KeyNOTWire_0[53]);
  xor XOR2_186 (KeyWire_0[116], N61, N707);
  xnor KeyGate_0_116(N739, keyIn_0_116, KeyWire_0[116]);
  xor XOR2_187 (KeyWire_0[117], N65, N708);
  xor KeyGate_0_117(KeyNOTWire_0[54], keyIn_0_117, KeyWire_0[117]);
  not KeyNOTGate_0_54(N740, KeyNOTWire_0[54]);
  xor XOR2_188 (KeyWire_0[118], N69, N709);
  xor KeyGate_0_118(KeyNOTWire_0[55], keyIn_0_118, KeyWire_0[118]);
  not KeyNOTGate_0_55(N741, KeyNOTWire_0[55]);
xor XOR2_189 (N742, N73, N710);
  xor XOR2_190 (KeyWire_0[119], N77, N711);
  xor KeyGate_0_119(N743, keyIn_0_119, KeyWire_0[119]);
  xor XOR2_191 (KeyWire_0[120], N81, N712);
  xor KeyGate_0_120(N744, keyIn_0_120, KeyWire_0[120]);
  xor XOR2_192 (KeyWire_0[121], N85, N713);
  xor KeyGate_0_121(KeyNOTWire_0[56], keyIn_0_121, KeyWire_0[121]);
  not KeyNOTGate_0_56(N745, KeyNOTWire_0[56]);
  xor XOR2_193 (KeyWire_0[122], N89, N714);
  xor KeyGate_0_122(N746, keyIn_0_122, KeyWire_0[122]);
xor XOR2_194 (N747, N93, N715);
xor XOR2_195 (N748, N97, N716);
xor XOR2_196 (N749, N101, N717);
  xor XOR2_197 (KeyWire_0[123], N105, N718);
  xor KeyGate_0_123(N750, keyIn_0_123, KeyWire_0[123]);
xor XOR2_198 (N751, N109, N719);
  xor XOR2_199 (KeyWire_0[124], N113, N720);
  xor KeyGate_0_124(KeyNOTWire_0[57], keyIn_0_124, KeyWire_0[124]);
  not KeyNOTGate_0_57(N752, KeyNOTWire_0[57]);
  xor XOR2_200 (KeyWire_0[125], N117, N721);
  xor KeyGate_0_125(KeyNOTWire_0[58], keyIn_0_125, KeyWire_0[125]);
  not KeyNOTGate_0_58(N753, KeyNOTWire_0[58]);
  xor XOR2_201 (KeyWire_0[126], N121, N722);
  xnor KeyGate_0_126(KeyNOTWire_0[59], keyIn_0_126, KeyWire_0[126]);
  not KeyNOTGate_0_59(N754, KeyNOTWire_0[59]);
  xor XOR2_202 (KeyWire_0[127], N125, N723);
  xor KeyGate_0_127(N755, keyIn_0_127, KeyWire_0[127]);

endmodule
